magic
tech scmos
timestamp 1681620392
<< metal1 >>
rect -10 -3 10 3
<< metal2 >>
rect -10 -3 10 3
<< gv1 >>
rect -9 -1 -7 1
rect -4 -1 -2 1
rect 1 -1 3 1
rect 6 -1 8 1
<< end >>
