magic
tech scmos
timestamp 1681620392
<< nwell >>
rect 20 740 280 1000
rect 15 604 286 652
rect 14 475 286 604
rect 14 425 285 475
rect 142 424 285 425
rect -6 253 303 338
rect -3 249 303 253
rect -3 11 11 249
rect 286 11 303 249
rect -3 -3 303 11
<< ntransistor >>
rect 19 353 21 383
rect 27 353 29 383
rect 44 353 46 383
rect 52 353 54 383
rect 60 353 62 383
rect 68 353 70 383
rect 76 353 78 383
rect 84 353 86 383
rect 92 353 94 383
rect 100 353 102 383
rect 108 353 110 383
rect 116 353 118 383
rect 124 353 126 383
rect 132 353 134 383
rect 140 353 142 383
rect 148 353 150 383
rect 198 353 200 383
rect 206 353 208 383
rect 214 353 216 383
rect 222 353 224 383
rect 230 353 232 383
rect 238 353 240 383
rect 246 353 248 383
rect 254 353 256 383
rect 262 353 264 383
rect 270 353 272 383
rect 278 353 280 383
rect 286 353 288 383
rect 38 216 138 219
rect 38 171 138 174
rect 38 150 138 153
rect 38 106 138 109
rect 38 85 138 88
rect 38 41 138 44
rect 162 216 262 219
rect 162 171 262 174
rect 162 150 262 153
rect 162 106 262 109
rect 162 85 262 88
rect 162 41 262 44
<< ptransistor >>
rect 38 624 138 627
rect 38 580 138 583
rect 38 559 138 562
rect 38 516 138 519
rect 38 495 138 498
rect 38 451 138 454
rect 162 624 262 627
rect 162 580 262 583
rect 162 559 262 562
rect 162 516 262 519
rect 162 495 262 498
rect 162 451 262 454
rect 19 269 21 321
rect 27 269 29 321
rect 44 269 46 321
rect 52 269 54 321
rect 60 269 62 321
rect 68 269 70 321
rect 76 269 78 321
rect 84 269 86 321
rect 92 269 94 321
rect 100 269 102 321
rect 108 269 110 321
rect 116 269 118 321
rect 124 269 126 321
rect 132 269 134 321
rect 140 269 142 321
rect 148 269 150 321
rect 198 269 200 321
rect 206 269 208 321
rect 214 269 216 321
rect 222 269 224 321
rect 230 269 232 321
rect 238 269 240 321
rect 246 269 248 321
rect 254 269 256 321
rect 262 269 264 321
rect 270 269 272 321
rect 278 269 280 321
rect 286 269 288 321
<< ndiffusion >>
rect 13 353 19 383
rect 21 353 27 383
rect 29 353 35 383
rect 38 353 44 383
rect 46 353 52 383
rect 54 353 60 383
rect 62 353 68 383
rect 70 353 76 383
rect 78 353 84 383
rect 86 353 92 383
rect 94 353 100 383
rect 102 353 108 383
rect 110 353 116 383
rect 118 353 124 383
rect 126 353 132 383
rect 134 353 140 383
rect 142 353 148 383
rect 150 353 156 383
rect 192 353 198 383
rect 200 353 206 383
rect 208 353 214 383
rect 216 353 222 383
rect 224 353 230 383
rect 232 353 238 383
rect 240 353 246 383
rect 248 353 254 383
rect 256 353 262 383
rect 264 353 270 383
rect 272 353 278 383
rect 280 353 286 383
rect 288 353 293 383
rect 47 350 50 353
rect 63 350 67 353
rect 79 350 83 353
rect 111 350 115 353
rect 192 350 197 353
rect 209 350 213 353
rect 225 350 228 353
rect 241 350 245 353
rect 257 350 261 353
rect 273 350 276 353
rect 289 350 293 353
rect 38 219 138 228
rect 38 174 138 216
rect 38 153 138 171
rect 38 109 138 150
rect 38 88 138 106
rect 38 44 138 85
rect 38 32 138 41
rect 38 31 43 32
rect 162 219 262 228
rect 162 174 262 216
rect 162 153 262 171
rect 162 109 262 150
rect 162 88 262 106
rect 162 44 262 85
rect 162 32 262 41
<< pdiffusion >>
rect 36 630 140 636
rect 160 630 264 636
rect 38 629 141 630
rect 159 629 262 630
rect 38 627 138 629
rect 38 583 138 624
rect 38 562 138 580
rect 38 519 138 559
rect 38 498 138 516
rect 38 454 138 495
rect 38 442 138 451
rect 162 627 262 629
rect 162 583 262 624
rect 162 562 262 580
rect 162 519 262 559
rect 162 498 262 516
rect 162 454 262 495
rect 162 442 262 451
rect 63 321 67 324
rect 79 321 83 324
rect 111 321 115 324
rect 192 321 197 324
rect 209 321 213 324
rect 225 321 228 324
rect 241 321 245 324
rect 257 321 261 324
rect 273 321 276 324
rect 289 321 293 324
rect 13 269 19 321
rect 21 269 27 321
rect 29 269 35 321
rect 38 269 44 321
rect 46 269 52 321
rect 54 269 60 321
rect 62 269 68 321
rect 70 269 76 321
rect 78 269 84 321
rect 86 269 92 321
rect 94 269 100 321
rect 102 269 108 321
rect 110 269 116 321
rect 118 269 124 321
rect 126 269 132 321
rect 134 269 140 321
rect 142 269 148 321
rect 150 269 156 321
rect 192 269 198 321
rect 200 269 206 321
rect 208 269 214 321
rect 216 269 222 321
rect 224 269 230 321
rect 232 269 238 321
rect 240 269 246 321
rect 248 269 254 321
rect 256 269 262 321
rect 264 269 270 321
rect 272 269 278 321
rect 280 269 286 321
rect 288 269 293 321
rect 79 266 83 269
rect 192 266 197 269
rect 241 266 245 269
rect 289 257 293 269
<< psubstratepdiff >>
rect 0 657 300 670
rect 0 420 11 657
rect 117 420 147 421
rect 153 420 183 421
rect 289 420 300 657
rect 0 410 300 420
rect 0 348 6 410
rect 0 345 7 348
rect 15 345 23 348
rect 47 347 50 350
rect 31 345 50 347
rect 63 347 67 350
rect 79 347 83 350
rect 63 345 84 347
rect 111 348 115 350
rect 97 345 135 348
rect 192 348 197 350
rect 209 348 213 350
rect 225 348 228 350
rect 148 345 228 348
rect 241 348 245 350
rect 257 348 261 350
rect 273 348 276 350
rect 241 345 276 348
rect 293 350 300 410
rect 289 345 300 350
rect 0 344 50 345
rect 63 344 300 345
rect 0 341 300 344
rect 14 230 281 246
rect 14 31 30 230
rect 38 228 138 230
rect 43 31 138 32
rect 14 30 138 31
rect 143 30 157 230
rect 162 228 262 230
rect 162 30 262 32
rect 270 30 281 230
rect 14 14 281 30
<< nsubstratendiff >>
rect 19 636 281 648
rect 19 630 36 636
rect 140 630 160 636
rect 264 630 281 636
rect 19 440 30 630
rect 141 629 159 630
rect 38 440 138 442
rect 142 440 158 629
rect 162 440 262 442
rect 270 440 281 630
rect 19 430 281 440
rect 0 329 300 332
rect 0 326 7 329
rect 0 261 6 326
rect 15 326 23 329
rect 31 326 50 329
rect 63 326 84 329
rect 63 324 67 326
rect 79 324 83 326
rect 97 326 122 329
rect 111 324 115 326
rect 135 326 228 329
rect 192 324 197 326
rect 209 324 213 326
rect 225 324 228 326
rect 241 326 276 329
rect 241 324 245 326
rect 257 324 261 326
rect 273 324 276 326
rect 289 324 300 329
rect 36 261 43 265
rect 79 265 83 266
rect 192 265 197 266
rect 241 265 245 266
rect 56 261 289 265
rect 0 257 289 261
rect 293 257 300 324
rect 0 252 300 257
rect 0 8 8 252
rect 289 8 300 252
rect 0 0 300 8
<< polysilicon >>
rect 6 714 21 717
rect 24 714 39 717
rect 12 702 15 714
rect 24 711 27 714
rect 36 711 39 714
rect 24 708 39 711
rect 24 702 27 708
rect 36 702 39 708
rect 42 714 45 717
rect 42 711 51 714
rect 42 702 45 711
rect 48 708 51 711
rect 54 708 57 717
rect 48 705 57 708
rect 54 702 57 705
rect 60 714 63 717
rect 60 711 69 714
rect 60 702 63 711
rect 66 708 69 711
rect 72 708 75 717
rect 66 705 75 708
rect 72 702 75 705
rect 78 714 93 717
rect 96 714 111 717
rect 78 711 81 714
rect 96 711 99 714
rect 108 711 111 714
rect 78 708 93 711
rect 96 708 111 711
rect 207 714 222 717
rect 78 705 81 708
rect 78 702 93 705
rect 96 702 99 708
rect 105 702 108 708
rect 207 702 210 714
rect 213 708 216 714
rect 219 702 222 714
rect 225 714 240 717
rect 225 705 228 714
rect 237 705 240 714
rect 243 714 258 717
rect 261 714 276 717
rect 279 714 294 717
rect 243 711 246 714
rect 243 708 258 711
rect 255 705 258 708
rect 267 705 270 714
rect 279 711 282 714
rect 279 708 294 711
rect 291 705 294 708
rect 225 702 240 705
rect 243 702 258 705
rect 261 702 276 705
rect 279 702 294 705
rect 54 689 69 692
rect 72 689 87 692
rect 90 689 105 692
rect 54 680 57 689
rect 72 686 75 689
rect 90 686 93 689
rect 72 683 87 686
rect 90 683 105 686
rect 72 680 75 683
rect 102 680 105 683
rect 54 677 69 680
rect 72 677 87 680
rect 90 677 105 680
rect 31 624 38 627
rect 138 624 141 627
rect 31 583 37 624
rect 139 583 141 624
rect 31 580 38 583
rect 138 580 141 583
rect 31 562 37 580
rect 139 562 141 580
rect 31 559 38 562
rect 138 559 141 562
rect 31 519 37 559
rect 139 519 141 559
rect 31 516 38 519
rect 138 516 141 519
rect 31 498 37 516
rect 139 498 141 516
rect 31 495 38 498
rect 138 495 141 498
rect 31 454 37 495
rect 139 454 141 495
rect 31 451 38 454
rect 138 451 141 454
rect 159 624 162 627
rect 262 624 269 627
rect 159 583 161 624
rect 263 583 269 624
rect 159 580 162 583
rect 262 580 269 583
rect 159 562 161 580
rect 263 562 269 580
rect 159 559 162 562
rect 262 559 269 562
rect 159 519 161 559
rect 263 519 269 559
rect 159 516 162 519
rect 262 516 269 519
rect 159 498 161 516
rect 263 498 269 516
rect 159 495 162 498
rect 262 495 269 498
rect 159 454 161 495
rect 263 454 269 495
rect 159 451 162 454
rect 262 451 269 454
rect 111 395 126 405
rect 191 395 210 405
rect 274 395 290 405
rect 193 390 208 395
rect 19 383 21 385
rect 24 384 35 390
rect 44 384 78 386
rect 27 383 29 384
rect 44 383 46 384
rect 52 383 54 384
rect 60 383 62 384
rect 68 383 70 384
rect 76 383 78 384
rect 84 384 118 386
rect 84 383 86 384
rect 92 383 94 384
rect 100 383 102 384
rect 108 383 110 384
rect 116 383 118 384
rect 124 383 126 385
rect 132 383 134 385
rect 140 383 142 385
rect 148 383 150 385
rect 198 383 200 390
rect 206 384 216 386
rect 206 383 208 384
rect 214 383 216 384
rect 222 384 232 386
rect 222 383 224 384
rect 230 383 232 384
rect 238 383 240 385
rect 246 383 248 385
rect 254 384 264 386
rect 254 383 256 384
rect 262 383 264 384
rect 270 384 280 386
rect 270 383 272 384
rect 278 383 280 384
rect 286 383 288 386
rect 19 352 21 353
rect 27 352 29 353
rect 8 350 21 352
rect 8 346 14 350
rect 24 346 30 352
rect 44 350 46 353
rect 52 351 54 353
rect 60 351 62 353
rect 51 345 62 351
rect 68 350 70 353
rect 76 350 78 353
rect 84 352 86 353
rect 92 352 94 353
rect 84 349 96 352
rect 100 350 102 353
rect 108 350 110 353
rect 116 350 118 353
rect 124 352 126 353
rect 132 352 134 353
rect 140 352 142 353
rect 148 352 150 353
rect 124 350 150 352
rect 198 352 200 353
rect 206 352 208 353
rect 198 350 208 352
rect 214 352 216 353
rect 222 352 224 353
rect 214 350 224 352
rect 230 352 232 353
rect 238 352 240 353
rect 85 346 96 349
rect 136 346 147 350
rect 229 346 240 352
rect 246 352 248 353
rect 254 352 256 353
rect 246 350 256 352
rect 262 352 264 353
rect 270 352 272 353
rect 262 350 272 352
rect 278 352 280 353
rect 286 352 288 353
rect 277 346 288 352
rect 31 334 147 340
rect 8 324 14 328
rect 8 322 21 324
rect 24 322 30 328
rect 19 321 21 322
rect 27 321 29 322
rect 44 321 46 323
rect 51 322 62 328
rect 52 321 54 322
rect 60 321 62 322
rect 85 324 96 328
rect 68 321 70 323
rect 76 321 78 323
rect 84 322 96 324
rect 84 321 86 322
rect 92 321 94 322
rect 100 321 102 323
rect 108 321 110 323
rect 123 324 134 328
rect 116 321 118 323
rect 123 322 150 324
rect 124 321 126 322
rect 132 321 134 322
rect 140 321 142 322
rect 148 321 150 322
rect 198 323 208 325
rect 198 321 200 323
rect 206 321 208 323
rect 214 323 224 325
rect 214 321 216 323
rect 222 321 224 323
rect 229 322 240 328
rect 230 321 232 322
rect 238 321 240 322
rect 246 322 256 324
rect 246 321 248 322
rect 254 321 256 322
rect 262 322 272 324
rect 262 321 264 322
rect 270 321 272 322
rect 277 322 288 328
rect 278 321 280 322
rect 286 321 288 322
rect 19 268 21 269
rect 27 268 29 269
rect 44 268 46 269
rect 52 268 54 269
rect 60 268 62 269
rect 68 268 70 269
rect 76 268 78 269
rect 10 262 21 268
rect 24 262 35 268
rect 44 266 78 268
rect 84 268 86 269
rect 92 268 94 269
rect 100 268 102 269
rect 108 268 110 269
rect 116 268 118 269
rect 84 266 118 268
rect 124 267 126 269
rect 132 267 134 269
rect 140 267 142 269
rect 148 267 150 269
rect 198 267 200 269
rect 206 268 208 269
rect 214 268 216 269
rect 206 266 216 268
rect 222 268 224 269
rect 230 268 232 269
rect 222 266 232 268
rect 238 267 240 269
rect 246 267 248 269
rect 254 268 256 269
rect 262 268 264 269
rect 254 266 264 268
rect 270 268 272 269
rect 278 268 280 269
rect 270 266 280 268
rect 286 267 288 269
rect 44 262 55 266
rect 31 216 38 219
rect 138 216 142 219
rect 31 174 37 216
rect 139 174 142 216
rect 31 171 38 174
rect 138 171 142 174
rect 31 153 37 171
rect 139 153 142 171
rect 31 150 38 153
rect 138 150 142 153
rect 31 109 37 150
rect 139 109 142 150
rect 31 106 38 109
rect 138 106 142 109
rect 31 88 37 106
rect 139 88 142 106
rect 31 85 38 88
rect 138 85 142 88
rect 31 44 37 85
rect 139 44 142 85
rect 31 41 38 44
rect 138 41 142 44
rect 158 216 162 219
rect 262 216 269 219
rect 158 174 161 216
rect 263 174 269 216
rect 158 171 162 174
rect 262 171 269 174
rect 158 153 161 171
rect 263 153 269 171
rect 158 150 162 153
rect 262 150 269 153
rect 158 109 161 150
rect 263 109 269 150
rect 158 106 162 109
rect 262 106 269 109
rect 158 88 161 106
rect 263 88 269 106
rect 158 85 162 88
rect 262 85 269 88
rect 158 44 161 85
rect 263 44 269 85
rect 158 41 162 44
rect 262 41 269 44
<< genericcontact >>
rect 2 664 4 666
rect 7 664 9 666
rect 12 664 14 666
rect 17 664 19 666
rect 22 664 24 666
rect 27 664 29 666
rect 32 664 34 666
rect 37 664 39 666
rect 42 664 44 666
rect 47 664 49 666
rect 52 664 54 666
rect 57 664 59 666
rect 62 664 64 666
rect 67 664 69 666
rect 72 664 74 666
rect 77 664 79 666
rect 82 664 84 666
rect 87 664 89 666
rect 92 664 94 666
rect 97 664 99 666
rect 102 664 104 666
rect 107 664 109 666
rect 112 664 114 666
rect 185 664 187 666
rect 190 664 192 666
rect 195 664 197 666
rect 200 664 202 666
rect 205 664 207 666
rect 210 664 212 666
rect 215 664 217 666
rect 220 664 222 666
rect 225 664 227 666
rect 230 664 232 666
rect 235 664 237 666
rect 240 664 242 666
rect 245 664 247 666
rect 250 664 252 666
rect 255 664 257 666
rect 260 664 262 666
rect 265 664 267 666
rect 270 664 272 666
rect 275 664 277 666
rect 280 664 282 666
rect 285 664 287 666
rect 290 664 292 666
rect 295 664 297 666
rect 2 659 4 661
rect 7 659 9 661
rect 12 659 14 661
rect 17 659 19 661
rect 22 659 24 661
rect 27 659 29 661
rect 32 659 34 661
rect 37 659 39 661
rect 42 659 44 661
rect 47 659 49 661
rect 52 659 54 661
rect 57 659 59 661
rect 62 659 64 661
rect 67 659 69 661
rect 72 659 74 661
rect 77 659 79 661
rect 82 659 84 661
rect 87 659 89 661
rect 92 659 94 661
rect 97 659 99 661
rect 102 659 104 661
rect 107 659 109 661
rect 112 659 114 661
rect 185 659 187 661
rect 190 659 192 661
rect 195 659 197 661
rect 200 659 202 661
rect 205 659 207 661
rect 210 659 212 661
rect 215 659 217 661
rect 220 659 222 661
rect 225 659 227 661
rect 230 659 232 661
rect 235 659 237 661
rect 240 659 242 661
rect 245 659 247 661
rect 250 659 252 661
rect 255 659 257 661
rect 260 659 262 661
rect 265 659 267 661
rect 270 659 272 661
rect 275 659 277 661
rect 280 659 282 661
rect 285 659 287 661
rect 290 659 292 661
rect 295 659 297 661
rect 291 653 293 655
rect 296 653 298 655
rect 2 651 4 653
rect 7 651 9 653
rect 291 648 293 650
rect 296 648 298 650
rect 2 646 4 648
rect 7 646 9 648
rect 149 644 151 646
rect 2 641 4 643
rect 7 641 9 643
rect 46 642 48 644
rect 51 642 53 644
rect 57 642 59 644
rect 67 642 69 644
rect 72 642 74 644
rect 82 642 84 644
rect 87 642 89 644
rect 97 642 99 644
rect 102 642 104 644
rect 112 642 114 644
rect 184 642 186 644
rect 194 642 196 644
rect 199 642 201 644
rect 209 642 211 644
rect 214 642 216 644
rect 224 642 226 644
rect 229 642 231 644
rect 239 642 241 644
rect 245 642 247 644
rect 250 642 252 644
rect 291 643 293 645
rect 296 643 298 645
rect 2 636 4 638
rect 7 636 9 638
rect 21 637 23 639
rect 26 637 28 639
rect 46 637 48 639
rect 51 637 53 639
rect 57 637 59 639
rect 67 637 69 639
rect 72 637 74 639
rect 82 637 84 639
rect 87 637 89 639
rect 97 637 99 639
rect 102 637 104 639
rect 112 637 114 639
rect 184 637 186 639
rect 194 637 196 639
rect 199 637 201 639
rect 209 637 211 639
rect 214 637 216 639
rect 224 637 226 639
rect 229 637 231 639
rect 239 637 241 639
rect 245 637 247 639
rect 250 637 252 639
rect 272 637 274 639
rect 277 637 279 639
rect 291 638 293 640
rect 296 638 298 640
rect 149 634 151 636
rect 2 631 4 633
rect 7 631 9 633
rect 21 632 23 634
rect 26 632 28 634
rect 46 631 48 633
rect 51 631 53 633
rect 57 631 59 633
rect 67 631 69 633
rect 72 631 74 633
rect 82 631 84 633
rect 87 631 89 633
rect 97 631 99 633
rect 102 631 104 633
rect 112 631 114 633
rect 184 631 186 633
rect 194 631 196 633
rect 199 631 201 633
rect 209 631 211 633
rect 214 631 216 633
rect 224 631 226 633
rect 229 631 231 633
rect 239 631 241 633
rect 245 631 247 633
rect 250 631 252 633
rect 272 632 274 634
rect 277 632 279 634
rect 291 633 293 635
rect 296 633 298 635
rect 149 629 151 631
rect 2 626 4 628
rect 7 626 9 628
rect 21 627 23 629
rect 26 627 28 629
rect 272 627 274 629
rect 277 627 279 629
rect 291 628 293 630
rect 296 628 298 630
rect 149 624 151 626
rect 291 623 293 625
rect 296 623 298 625
rect 2 621 4 623
rect 7 621 9 623
rect 2 616 4 618
rect 7 616 9 618
rect 21 617 23 619
rect 26 617 28 619
rect 272 617 274 619
rect 277 617 279 619
rect 291 618 293 620
rect 296 618 298 620
rect 149 614 151 616
rect 2 611 4 613
rect 7 611 9 613
rect 21 612 23 614
rect 26 612 28 614
rect 33 611 35 613
rect 272 612 274 614
rect 277 612 279 614
rect 291 613 293 615
rect 296 613 298 615
rect 149 609 151 611
rect 265 609 267 611
rect 2 606 4 608
rect 7 606 9 608
rect 21 607 23 609
rect 26 607 28 609
rect 33 606 35 608
rect 272 607 274 609
rect 277 607 279 609
rect 291 608 293 610
rect 296 608 298 610
rect 57 605 59 607
rect 62 605 64 607
rect 67 605 69 607
rect 72 605 74 607
rect 77 605 79 607
rect 82 605 84 607
rect 87 605 89 607
rect 92 605 94 607
rect 97 605 99 607
rect 102 605 104 607
rect 107 605 109 607
rect 112 605 114 607
rect 117 605 119 607
rect 149 604 151 606
rect 181 605 183 607
rect 186 605 188 607
rect 191 605 193 607
rect 196 605 198 607
rect 201 605 203 607
rect 206 605 208 607
rect 211 605 213 607
rect 216 605 218 607
rect 221 605 223 607
rect 226 605 228 607
rect 231 605 233 607
rect 236 605 238 607
rect 241 605 243 607
rect 265 604 267 606
rect 291 603 293 605
rect 296 603 298 605
rect 2 601 4 603
rect 7 601 9 603
rect 33 601 35 603
rect 57 600 59 602
rect 62 600 64 602
rect 67 600 69 602
rect 72 600 74 602
rect 77 600 79 602
rect 82 600 84 602
rect 87 600 89 602
rect 92 600 94 602
rect 97 600 99 602
rect 102 600 104 602
rect 107 600 109 602
rect 112 600 114 602
rect 117 600 119 602
rect 181 600 183 602
rect 186 600 188 602
rect 191 600 193 602
rect 196 600 198 602
rect 201 600 203 602
rect 206 600 208 602
rect 211 600 213 602
rect 216 600 218 602
rect 221 600 223 602
rect 226 600 228 602
rect 231 600 233 602
rect 236 600 238 602
rect 241 600 243 602
rect 265 599 267 601
rect 2 596 4 598
rect 7 596 9 598
rect 21 597 23 599
rect 26 597 28 599
rect 33 596 35 598
rect 272 597 274 599
rect 277 597 279 599
rect 291 598 293 600
rect 296 598 298 600
rect 149 594 151 596
rect 265 594 267 596
rect 2 591 4 593
rect 7 591 9 593
rect 21 592 23 594
rect 26 592 28 594
rect 272 592 274 594
rect 277 592 279 594
rect 291 593 293 595
rect 296 593 298 595
rect 149 589 151 591
rect 2 586 4 588
rect 7 586 9 588
rect 21 587 23 589
rect 26 587 28 589
rect 272 587 274 589
rect 277 587 279 589
rect 291 588 293 590
rect 296 588 298 590
rect 149 584 151 586
rect 291 583 293 585
rect 296 583 298 585
rect 2 581 4 583
rect 7 581 9 583
rect 2 576 4 578
rect 7 576 9 578
rect 21 577 23 579
rect 26 577 28 579
rect 272 577 274 579
rect 277 577 279 579
rect 291 578 293 580
rect 296 578 298 580
rect 2 571 4 573
rect 7 571 9 573
rect 21 572 23 574
rect 26 572 28 574
rect 62 573 64 575
rect 67 573 69 575
rect 77 573 79 575
rect 82 573 84 575
rect 92 573 94 575
rect 97 573 99 575
rect 107 573 109 575
rect 112 573 114 575
rect 149 574 151 576
rect 185 573 187 575
rect 190 573 192 575
rect 200 573 202 575
rect 205 573 207 575
rect 215 573 217 575
rect 220 573 222 575
rect 230 573 232 575
rect 235 573 237 575
rect 272 572 274 574
rect 277 572 279 574
rect 291 573 293 575
rect 296 573 298 575
rect 149 569 151 571
rect 2 566 4 568
rect 7 566 9 568
rect 21 567 23 569
rect 26 567 28 569
rect 62 567 64 569
rect 67 567 69 569
rect 77 567 79 569
rect 82 567 84 569
rect 92 567 94 569
rect 97 567 99 569
rect 107 567 109 569
rect 112 567 114 569
rect 185 567 187 569
rect 190 567 192 569
rect 200 567 202 569
rect 205 567 207 569
rect 215 567 217 569
rect 220 567 222 569
rect 230 567 232 569
rect 235 567 237 569
rect 272 567 274 569
rect 277 567 279 569
rect 291 568 293 570
rect 296 568 298 570
rect 149 564 151 566
rect 291 563 293 565
rect 296 563 298 565
rect 2 561 4 563
rect 7 561 9 563
rect 2 556 4 558
rect 7 556 9 558
rect 21 557 23 559
rect 26 557 28 559
rect 272 557 274 559
rect 277 557 279 559
rect 291 558 293 560
rect 296 558 298 560
rect 149 554 151 556
rect 2 551 4 553
rect 7 551 9 553
rect 21 552 23 554
rect 26 552 28 554
rect 272 552 274 554
rect 277 552 279 554
rect 291 553 293 555
rect 296 553 298 555
rect 149 549 151 551
rect 2 546 4 548
rect 7 546 9 548
rect 21 547 23 549
rect 26 547 28 549
rect 33 546 35 548
rect 265 546 267 548
rect 272 547 274 549
rect 277 547 279 549
rect 291 548 293 550
rect 296 548 298 550
rect 149 544 151 546
rect 291 543 293 545
rect 296 543 298 545
rect 2 541 4 543
rect 7 541 9 543
rect 33 541 35 543
rect 57 540 59 542
rect 62 540 64 542
rect 67 540 69 542
rect 72 540 74 542
rect 77 540 79 542
rect 82 540 84 542
rect 87 540 89 542
rect 92 540 94 542
rect 97 540 99 542
rect 102 540 104 542
rect 107 540 109 542
rect 112 540 114 542
rect 117 540 119 542
rect 181 540 183 542
rect 186 540 188 542
rect 191 540 193 542
rect 196 540 198 542
rect 201 540 203 542
rect 206 540 208 542
rect 211 540 213 542
rect 216 540 218 542
rect 221 540 223 542
rect 226 540 228 542
rect 231 540 233 542
rect 236 540 238 542
rect 241 540 243 542
rect 265 541 267 543
rect 2 536 4 538
rect 7 536 9 538
rect 21 537 23 539
rect 26 537 28 539
rect 33 536 35 538
rect 57 535 59 537
rect 62 535 64 537
rect 67 535 69 537
rect 72 535 74 537
rect 77 535 79 537
rect 82 535 84 537
rect 87 535 89 537
rect 92 535 94 537
rect 97 535 99 537
rect 102 535 104 537
rect 107 535 109 537
rect 112 535 114 537
rect 117 535 119 537
rect 149 534 151 536
rect 181 535 183 537
rect 186 535 188 537
rect 191 535 193 537
rect 196 535 198 537
rect 201 535 203 537
rect 206 535 208 537
rect 211 535 213 537
rect 216 535 218 537
rect 221 535 223 537
rect 226 535 228 537
rect 231 535 233 537
rect 236 535 238 537
rect 241 535 243 537
rect 265 536 267 538
rect 272 537 274 539
rect 277 537 279 539
rect 291 538 293 540
rect 296 538 298 540
rect 2 531 4 533
rect 7 531 9 533
rect 21 532 23 534
rect 26 532 28 534
rect 33 531 35 533
rect 265 531 267 533
rect 272 532 274 534
rect 277 532 279 534
rect 291 533 293 535
rect 296 533 298 535
rect 149 529 151 531
rect 2 526 4 528
rect 7 526 9 528
rect 21 527 23 529
rect 26 527 28 529
rect 272 527 274 529
rect 277 527 279 529
rect 291 528 293 530
rect 296 528 298 530
rect 149 524 151 526
rect 291 523 293 525
rect 296 523 298 525
rect 2 521 4 523
rect 7 521 9 523
rect 2 516 4 518
rect 7 516 9 518
rect 21 517 23 519
rect 26 517 28 519
rect 272 517 274 519
rect 277 517 279 519
rect 291 518 293 520
rect 296 518 298 520
rect 149 514 151 516
rect 2 511 4 513
rect 7 511 9 513
rect 21 512 23 514
rect 26 512 28 514
rect 272 512 274 514
rect 277 512 279 514
rect 291 513 293 515
rect 296 513 298 515
rect 62 509 64 511
rect 67 509 69 511
rect 77 509 79 511
rect 82 509 84 511
rect 92 509 94 511
rect 97 509 99 511
rect 107 509 109 511
rect 112 509 114 511
rect 149 509 151 511
rect 184 509 186 511
rect 189 509 191 511
rect 199 509 201 511
rect 204 509 206 511
rect 214 509 216 511
rect 219 509 221 511
rect 229 509 231 511
rect 234 509 236 511
rect 2 506 4 508
rect 7 506 9 508
rect 21 507 23 509
rect 26 507 28 509
rect 272 507 274 509
rect 277 507 279 509
rect 291 508 293 510
rect 296 508 298 510
rect 62 503 64 505
rect 67 503 69 505
rect 77 503 79 505
rect 82 503 84 505
rect 92 503 94 505
rect 97 503 99 505
rect 107 503 109 505
rect 112 503 114 505
rect 149 504 151 506
rect 184 503 186 505
rect 189 503 191 505
rect 199 503 201 505
rect 204 503 206 505
rect 214 503 216 505
rect 219 503 221 505
rect 229 503 231 505
rect 234 503 236 505
rect 291 503 293 505
rect 296 503 298 505
rect 2 501 4 503
rect 7 501 9 503
rect 2 496 4 498
rect 7 496 9 498
rect 21 497 23 499
rect 26 497 28 499
rect 272 497 274 499
rect 277 497 279 499
rect 291 498 293 500
rect 296 498 298 500
rect 149 494 151 496
rect 2 491 4 493
rect 7 491 9 493
rect 21 492 23 494
rect 26 492 28 494
rect 272 492 274 494
rect 277 492 279 494
rect 291 493 293 495
rect 296 493 298 495
rect 149 489 151 491
rect 2 486 4 488
rect 7 486 9 488
rect 21 487 23 489
rect 26 487 28 489
rect 272 487 274 489
rect 277 487 279 489
rect 291 488 293 490
rect 296 488 298 490
rect 149 484 151 486
rect 291 483 293 485
rect 296 483 298 485
rect 2 481 4 483
rect 7 481 9 483
rect 265 481 267 483
rect 2 476 4 478
rect 7 476 9 478
rect 21 477 23 479
rect 26 477 28 479
rect 33 478 35 480
rect 57 476 59 478
rect 62 476 64 478
rect 67 476 69 478
rect 72 476 74 478
rect 77 476 79 478
rect 82 476 84 478
rect 87 476 89 478
rect 92 476 94 478
rect 97 476 99 478
rect 102 476 104 478
rect 107 476 109 478
rect 112 476 114 478
rect 117 476 119 478
rect 181 476 183 478
rect 186 476 188 478
rect 191 476 193 478
rect 196 476 198 478
rect 201 476 203 478
rect 206 476 208 478
rect 211 476 213 478
rect 216 476 218 478
rect 221 476 223 478
rect 226 476 228 478
rect 231 476 233 478
rect 236 476 238 478
rect 241 476 243 478
rect 265 476 267 478
rect 272 477 274 479
rect 277 477 279 479
rect 291 478 293 480
rect 296 478 298 480
rect 2 471 4 473
rect 7 471 9 473
rect 21 472 23 474
rect 26 472 28 474
rect 33 473 35 475
rect 149 474 151 476
rect 57 471 59 473
rect 62 471 64 473
rect 67 471 69 473
rect 72 471 74 473
rect 77 471 79 473
rect 82 471 84 473
rect 87 471 89 473
rect 92 471 94 473
rect 97 471 99 473
rect 102 471 104 473
rect 107 471 109 473
rect 112 471 114 473
rect 117 471 119 473
rect 181 471 183 473
rect 186 471 188 473
rect 191 471 193 473
rect 196 471 198 473
rect 201 471 203 473
rect 206 471 208 473
rect 211 471 213 473
rect 216 471 218 473
rect 221 471 223 473
rect 226 471 228 473
rect 231 471 233 473
rect 236 471 238 473
rect 241 471 243 473
rect 265 471 267 473
rect 272 472 274 474
rect 277 472 279 474
rect 291 473 293 475
rect 296 473 298 475
rect 2 466 4 468
rect 7 466 9 468
rect 21 467 23 469
rect 26 467 28 469
rect 33 468 35 470
rect 149 469 151 471
rect 265 466 267 468
rect 272 467 274 469
rect 277 467 279 469
rect 291 468 293 470
rect 296 468 298 470
rect 33 463 35 465
rect 149 464 151 466
rect 291 463 293 465
rect 296 463 298 465
rect 2 461 4 463
rect 7 461 9 463
rect 265 461 267 463
rect 2 456 4 458
rect 7 456 9 458
rect 21 457 23 459
rect 26 457 28 459
rect 33 458 35 460
rect 265 456 267 458
rect 272 457 274 459
rect 277 457 279 459
rect 291 458 293 460
rect 296 458 298 460
rect 2 451 4 453
rect 7 451 9 453
rect 21 452 23 454
rect 26 452 28 454
rect 33 453 35 455
rect 149 454 151 456
rect 272 452 274 454
rect 277 452 279 454
rect 291 453 293 455
rect 296 453 298 455
rect 149 449 151 451
rect 2 446 4 448
rect 7 446 9 448
rect 21 447 23 449
rect 26 447 28 449
rect 272 447 274 449
rect 277 447 279 449
rect 291 448 293 450
rect 296 448 298 450
rect 62 444 64 446
rect 67 444 69 446
rect 77 444 79 446
rect 82 444 84 446
rect 92 444 94 446
rect 97 444 99 446
rect 107 444 109 446
rect 112 444 114 446
rect 149 444 151 446
rect 185 444 187 446
rect 190 444 192 446
rect 200 444 202 446
rect 205 444 207 446
rect 215 444 217 446
rect 220 444 222 446
rect 230 444 232 446
rect 235 444 237 446
rect 291 443 293 445
rect 296 443 298 445
rect 2 441 4 443
rect 7 441 9 443
rect 2 436 4 438
rect 7 436 9 438
rect 21 437 23 439
rect 26 437 28 439
rect 52 438 54 440
rect 62 438 64 440
rect 67 438 69 440
rect 77 438 79 440
rect 82 438 84 440
rect 92 438 94 440
rect 97 438 99 440
rect 107 438 109 440
rect 112 438 114 440
rect 185 438 187 440
rect 190 438 192 440
rect 200 438 202 440
rect 205 438 207 440
rect 215 438 217 440
rect 220 438 222 440
rect 230 438 232 440
rect 235 438 237 440
rect 245 438 247 440
rect 272 437 274 439
rect 277 437 279 439
rect 291 438 293 440
rect 296 438 298 440
rect 149 434 151 436
rect 2 431 4 433
rect 7 431 9 433
rect 21 432 23 434
rect 26 432 28 434
rect 47 432 49 434
rect 52 432 54 434
rect 57 432 59 434
rect 62 432 64 434
rect 67 432 69 434
rect 72 432 74 434
rect 77 432 79 434
rect 82 432 84 434
rect 87 432 89 434
rect 92 432 94 434
rect 97 432 99 434
rect 102 432 104 434
rect 107 432 109 434
rect 112 432 114 434
rect 185 432 187 434
rect 190 432 192 434
rect 195 432 197 434
rect 200 432 202 434
rect 205 432 207 434
rect 210 432 212 434
rect 215 432 217 434
rect 220 432 222 434
rect 225 432 227 434
rect 230 432 232 434
rect 235 432 237 434
rect 240 432 242 434
rect 245 432 247 434
rect 250 432 252 434
rect 272 432 274 434
rect 277 432 279 434
rect 291 433 293 435
rect 296 433 298 435
rect 291 428 293 430
rect 296 428 298 430
rect 2 426 4 428
rect 7 426 9 428
rect 291 423 293 425
rect 296 423 298 425
rect 2 421 4 423
rect 7 421 9 423
rect 291 418 293 420
rect 296 418 298 420
rect 2 416 4 418
rect 7 416 9 418
rect 16 416 18 418
rect 21 416 23 418
rect 26 416 28 418
rect 40 416 42 418
rect 45 416 47 418
rect 50 416 52 418
rect 55 416 57 418
rect 60 416 62 418
rect 65 416 67 418
rect 70 416 72 418
rect 75 416 77 418
rect 80 416 82 418
rect 85 416 87 418
rect 90 416 92 418
rect 95 416 97 418
rect 100 416 102 418
rect 105 416 107 418
rect 110 416 112 418
rect 149 416 151 418
rect 185 416 187 418
rect 190 416 192 418
rect 195 416 197 418
rect 200 416 202 418
rect 205 416 207 418
rect 210 416 212 418
rect 215 416 217 418
rect 220 416 222 418
rect 225 416 227 418
rect 230 416 232 418
rect 235 416 237 418
rect 240 416 242 418
rect 245 416 247 418
rect 250 416 252 418
rect 255 416 257 418
rect 260 416 262 418
rect 265 416 267 418
rect 270 416 272 418
rect 275 416 277 418
rect 280 416 282 418
rect 285 416 287 418
rect 291 413 293 415
rect 296 413 298 415
rect 16 411 18 413
rect 21 411 23 413
rect 26 411 28 413
rect 40 411 42 413
rect 45 411 47 413
rect 50 411 52 413
rect 55 411 57 413
rect 60 411 62 413
rect 65 411 67 413
rect 70 411 72 413
rect 75 411 77 413
rect 80 411 82 413
rect 85 411 87 413
rect 90 411 92 413
rect 95 411 97 413
rect 100 411 102 413
rect 105 411 107 413
rect 110 411 112 413
rect 149 411 151 413
rect 185 411 187 413
rect 190 411 192 413
rect 195 411 197 413
rect 200 411 202 413
rect 205 411 207 413
rect 210 411 212 413
rect 215 411 217 413
rect 220 411 222 413
rect 225 411 227 413
rect 230 411 232 413
rect 235 411 237 413
rect 240 411 242 413
rect 245 411 247 413
rect 250 411 252 413
rect 255 411 257 413
rect 260 411 262 413
rect 265 411 267 413
rect 270 411 272 413
rect 275 411 277 413
rect 280 411 282 413
rect 285 411 287 413
rect 2 404 4 406
rect 296 403 298 405
rect 112 401 114 403
rect 117 401 119 403
rect 122 401 124 403
rect 276 401 278 403
rect 281 401 283 403
rect 286 401 288 403
rect 2 399 4 401
rect 112 396 114 398
rect 117 396 119 398
rect 122 396 124 398
rect 194 396 196 398
rect 199 396 201 398
rect 204 396 206 398
rect 276 396 278 398
rect 281 396 283 398
rect 286 396 288 398
rect 2 394 4 396
rect 296 393 298 395
rect 194 391 196 393
rect 199 391 201 393
rect 204 391 206 393
rect 2 389 4 391
rect 26 386 28 388
rect 31 386 33 388
rect 2 384 4 386
rect 296 383 298 385
rect 2 379 4 381
rect 152 379 154 381
rect 15 377 17 379
rect 23 377 25 379
rect 31 376 33 378
rect 40 376 42 378
rect 2 374 4 376
rect 48 375 50 377
rect 56 376 58 378
rect 64 375 66 377
rect 72 376 74 378
rect 80 375 82 377
rect 88 376 90 378
rect 104 377 106 379
rect 96 375 98 377
rect 112 375 114 377
rect 120 376 122 378
rect 128 375 130 377
rect 136 376 138 378
rect 144 376 146 378
rect 194 377 196 379
rect 202 377 204 379
rect 218 377 220 379
rect 226 377 228 379
rect 234 377 236 379
rect 242 377 244 379
rect 250 377 252 379
rect 258 377 260 379
rect 266 377 268 379
rect 274 377 276 379
rect 282 377 284 379
rect 290 377 292 379
rect 152 374 154 376
rect 15 372 17 374
rect 31 371 33 373
rect 40 371 42 373
rect 56 371 58 373
rect 72 371 74 373
rect 88 371 90 373
rect 104 372 106 374
rect 120 371 122 373
rect 2 369 4 371
rect 128 370 130 372
rect 136 371 138 373
rect 144 371 146 373
rect 202 372 204 374
rect 210 371 212 373
rect 218 372 220 374
rect 234 372 236 374
rect 250 372 252 374
rect 266 372 268 374
rect 282 372 284 374
rect 296 373 298 375
rect 152 369 154 371
rect 15 367 17 369
rect 23 367 25 369
rect 31 366 33 368
rect 40 366 42 368
rect 2 364 4 366
rect 48 365 50 367
rect 56 366 58 368
rect 64 365 66 367
rect 72 366 74 368
rect 80 365 82 367
rect 88 366 90 368
rect 104 367 106 369
rect 96 365 98 367
rect 112 365 114 367
rect 120 366 122 368
rect 128 365 130 367
rect 136 366 138 368
rect 144 366 146 368
rect 194 367 196 369
rect 202 367 204 369
rect 210 366 212 368
rect 218 367 220 369
rect 226 367 228 369
rect 234 367 236 369
rect 242 367 244 369
rect 250 367 252 369
rect 258 367 260 369
rect 266 367 268 369
rect 274 367 276 369
rect 282 367 284 369
rect 290 367 292 369
rect 152 364 154 366
rect 15 362 17 364
rect 31 361 33 363
rect 40 361 42 363
rect 56 361 58 363
rect 72 361 74 363
rect 88 361 90 363
rect 104 362 106 364
rect 2 359 4 361
rect 128 360 130 362
rect 144 361 146 363
rect 202 362 204 364
rect 218 362 220 364
rect 234 362 236 364
rect 250 362 252 364
rect 266 362 268 364
rect 282 362 284 364
rect 296 363 298 365
rect 152 359 154 361
rect 23 357 25 359
rect 31 356 33 358
rect 2 354 4 356
rect 48 355 50 357
rect 56 356 58 358
rect 64 355 66 357
rect 72 356 74 358
rect 80 355 82 357
rect 88 356 90 358
rect 104 357 106 359
rect 96 355 98 357
rect 112 355 114 357
rect 128 355 130 357
rect 136 356 138 358
rect 194 357 196 359
rect 202 357 204 359
rect 218 357 220 359
rect 226 357 228 359
rect 234 357 236 359
rect 242 357 244 359
rect 250 357 252 359
rect 258 357 260 359
rect 266 357 268 359
rect 274 357 276 359
rect 282 357 284 359
rect 290 357 292 359
rect 152 354 154 356
rect 210 355 212 357
rect 296 353 298 355
rect 2 349 4 351
rect 10 348 12 350
rect 26 348 28 350
rect 53 347 55 349
rect 58 347 60 349
rect 87 348 89 350
rect 92 348 94 350
rect 138 348 140 350
rect 143 348 145 350
rect 231 348 233 350
rect 236 348 238 350
rect 279 348 281 350
rect 284 348 286 350
rect 2 344 4 346
rect 18 344 20 346
rect 39 343 41 345
rect 46 343 48 345
rect 65 343 67 345
rect 70 343 72 345
rect 75 343 77 345
rect 80 343 82 345
rect 100 344 102 346
rect 109 344 111 346
rect 125 344 127 346
rect 195 343 197 345
rect 200 343 202 345
rect 205 343 207 345
rect 210 343 212 345
rect 224 344 226 346
rect 243 343 245 345
rect 248 343 250 345
rect 258 343 260 345
rect 272 343 274 345
rect 291 343 293 345
rect 296 343 298 345
rect 33 336 35 338
rect 38 336 40 338
rect 81 336 83 338
rect 86 336 88 338
rect 138 336 140 338
rect 143 336 145 338
rect 3 328 5 330
rect 18 328 20 330
rect 39 328 41 330
rect 46 328 48 330
rect 65 328 67 330
rect 75 328 77 330
rect 80 328 82 330
rect 99 328 101 330
rect 110 328 112 330
rect 138 328 140 330
rect 195 328 197 330
rect 200 328 202 330
rect 210 328 212 330
rect 224 328 226 330
rect 243 328 245 330
rect 248 328 250 330
rect 258 328 260 330
rect 272 328 274 330
rect 296 329 298 331
rect 3 323 5 325
rect 10 324 12 326
rect 26 324 28 326
rect 53 324 55 326
rect 58 324 60 326
rect 87 324 89 326
rect 92 324 94 326
rect 125 324 127 326
rect 130 324 132 326
rect 231 324 233 326
rect 236 324 238 326
rect 279 324 281 326
rect 284 324 286 326
rect 296 324 298 326
rect 3 318 5 320
rect 23 317 25 319
rect 31 316 33 318
rect 48 317 50 319
rect 56 316 58 318
rect 72 316 74 318
rect 88 317 90 319
rect 104 316 106 318
rect 112 317 114 319
rect 120 317 122 319
rect 136 317 138 319
rect 144 317 146 319
rect 3 313 5 315
rect 64 313 66 315
rect 80 313 82 315
rect 15 311 17 313
rect 31 311 33 313
rect 40 311 42 313
rect 56 311 58 313
rect 72 311 74 313
rect 88 312 90 314
rect 96 313 98 315
rect 104 311 106 313
rect 120 312 122 314
rect 144 312 146 314
rect 194 313 196 315
rect 202 313 204 315
rect 210 313 212 315
rect 218 313 220 315
rect 226 313 228 315
rect 234 313 236 315
rect 242 313 244 315
rect 250 313 252 315
rect 258 313 260 315
rect 266 313 268 315
rect 274 313 276 315
rect 282 313 284 315
rect 290 313 292 315
rect 3 308 5 310
rect 15 306 17 308
rect 23 307 25 309
rect 31 306 33 308
rect 40 306 42 308
rect 48 307 50 309
rect 56 306 58 308
rect 72 306 74 308
rect 88 307 90 309
rect 104 306 106 308
rect 112 307 114 309
rect 120 307 122 309
rect 128 308 130 310
rect 144 307 146 309
rect 202 308 204 310
rect 218 308 220 310
rect 234 308 236 310
rect 250 308 252 310
rect 266 308 268 310
rect 282 308 284 310
rect 290 308 292 310
rect 152 306 154 308
rect 3 303 5 305
rect 64 303 66 305
rect 80 303 82 305
rect 15 301 17 303
rect 31 301 33 303
rect 40 301 42 303
rect 56 301 58 303
rect 72 301 74 303
rect 88 302 90 304
rect 96 303 98 305
rect 104 301 106 303
rect 120 302 122 304
rect 128 303 130 305
rect 136 304 138 306
rect 144 302 146 304
rect 194 303 196 305
rect 202 303 204 305
rect 210 303 212 305
rect 218 303 220 305
rect 226 303 228 305
rect 234 303 236 305
rect 242 303 244 305
rect 250 303 252 305
rect 258 303 260 305
rect 266 303 268 305
rect 274 303 276 305
rect 282 303 284 305
rect 290 303 292 305
rect 152 301 154 303
rect 3 298 5 300
rect 15 296 17 298
rect 23 297 25 299
rect 31 296 33 298
rect 40 296 42 298
rect 48 297 50 299
rect 56 296 58 298
rect 72 296 74 298
rect 88 297 90 299
rect 104 296 106 298
rect 112 297 114 299
rect 120 297 122 299
rect 128 298 130 300
rect 136 299 138 301
rect 144 297 146 299
rect 202 298 204 300
rect 218 298 220 300
rect 234 298 236 300
rect 250 298 252 300
rect 266 298 268 300
rect 282 298 284 300
rect 290 298 292 300
rect 152 296 154 298
rect 3 293 5 295
rect 64 293 66 295
rect 80 293 82 295
rect 15 291 17 293
rect 31 291 33 293
rect 40 291 42 293
rect 56 291 58 293
rect 72 291 74 293
rect 88 292 90 294
rect 96 293 98 295
rect 104 291 106 293
rect 120 292 122 294
rect 128 293 130 295
rect 136 294 138 296
rect 144 292 146 294
rect 202 293 204 295
rect 218 293 220 295
rect 234 293 236 295
rect 250 293 252 295
rect 266 293 268 295
rect 282 293 284 295
rect 290 293 292 295
rect 152 291 154 293
rect 3 288 5 290
rect 15 286 17 288
rect 23 287 25 289
rect 31 286 33 288
rect 40 286 42 288
rect 48 287 50 289
rect 56 286 58 288
rect 72 286 74 288
rect 88 287 90 289
rect 104 286 106 288
rect 112 287 114 289
rect 120 287 122 289
rect 128 288 130 290
rect 136 289 138 291
rect 144 287 146 289
rect 194 288 196 290
rect 202 288 204 290
rect 210 288 212 290
rect 218 288 220 290
rect 226 288 228 290
rect 234 288 236 290
rect 242 288 244 290
rect 250 288 252 290
rect 258 288 260 290
rect 266 288 268 290
rect 274 288 276 290
rect 282 288 284 290
rect 290 288 292 290
rect 152 286 154 288
rect 3 283 5 285
rect 64 283 66 285
rect 80 283 82 285
rect 15 281 17 283
rect 31 281 33 283
rect 40 281 42 283
rect 56 281 58 283
rect 72 281 74 283
rect 88 282 90 284
rect 96 283 98 285
rect 104 281 106 283
rect 120 282 122 284
rect 128 283 130 285
rect 136 284 138 286
rect 144 282 146 284
rect 194 283 196 285
rect 202 283 204 285
rect 210 283 212 285
rect 218 283 220 285
rect 226 283 228 285
rect 234 283 236 285
rect 242 283 244 285
rect 250 283 252 285
rect 258 283 260 285
rect 266 283 268 285
rect 274 283 276 285
rect 282 283 284 285
rect 290 283 292 285
rect 152 281 154 283
rect 3 278 5 280
rect 15 276 17 278
rect 23 277 25 279
rect 31 276 33 278
rect 40 276 42 278
rect 48 277 50 279
rect 56 276 58 278
rect 72 276 74 278
rect 88 277 90 279
rect 104 276 106 278
rect 112 277 114 279
rect 120 277 122 279
rect 128 278 130 280
rect 136 279 138 281
rect 144 277 146 279
rect 202 278 204 280
rect 218 278 220 280
rect 234 278 236 280
rect 250 278 252 280
rect 266 278 268 280
rect 282 278 284 280
rect 290 278 292 280
rect 152 276 154 278
rect 3 273 5 275
rect 64 273 66 275
rect 80 273 82 275
rect 15 271 17 273
rect 31 271 33 273
rect 40 271 42 273
rect 56 271 58 273
rect 72 271 74 273
rect 88 272 90 274
rect 96 273 98 275
rect 104 271 106 273
rect 120 272 122 274
rect 128 273 130 275
rect 144 272 146 274
rect 194 273 196 275
rect 202 273 204 275
rect 210 273 212 275
rect 218 273 220 275
rect 226 273 228 275
rect 234 273 236 275
rect 242 273 244 275
rect 250 273 252 275
rect 258 273 260 275
rect 266 273 268 275
rect 274 273 276 275
rect 282 273 284 275
rect 290 273 292 275
rect 152 271 154 273
rect 3 268 5 270
rect 290 268 292 270
rect 3 263 5 265
rect 12 264 14 266
rect 17 264 19 266
rect 26 264 28 266
rect 31 264 33 266
rect 46 264 48 266
rect 51 264 53 266
rect 60 260 62 262
rect 65 260 67 262
rect 70 260 72 262
rect 75 260 77 262
rect 80 260 82 262
rect 85 260 87 262
rect 90 260 92 262
rect 95 260 97 262
rect 100 260 102 262
rect 105 260 107 262
rect 110 260 112 262
rect 194 261 196 263
rect 242 262 244 264
rect 290 263 292 265
rect 3 258 5 260
rect 18 255 20 257
rect 23 255 25 257
rect 28 255 30 257
rect 33 255 35 257
rect 3 253 5 255
rect 55 254 57 256
rect 60 254 62 256
rect 65 254 67 256
rect 70 254 72 256
rect 75 254 77 256
rect 80 254 82 256
rect 85 254 87 256
rect 90 254 92 256
rect 95 254 97 256
rect 100 254 102 256
rect 105 254 107 256
rect 195 255 197 257
rect 200 255 202 257
rect 205 255 207 257
rect 210 255 212 257
rect 215 255 217 257
rect 220 255 222 257
rect 225 255 227 257
rect 241 256 243 258
rect 246 256 248 258
rect 251 256 253 258
rect 264 257 266 259
rect 269 257 271 259
rect 274 257 276 259
rect 279 257 281 259
rect 284 257 286 259
rect 290 258 292 260
rect 3 248 5 250
rect 291 248 293 250
rect 296 248 298 250
rect 3 243 5 245
rect 291 243 293 245
rect 296 243 298 245
rect 271 240 273 242
rect 277 240 279 242
rect 3 238 5 240
rect 18 237 20 239
rect 23 237 25 239
rect 28 237 30 239
rect 33 237 35 239
rect 54 238 56 240
rect 59 238 61 240
rect 64 238 66 240
rect 69 238 71 240
rect 74 238 76 240
rect 79 238 81 240
rect 84 238 86 240
rect 89 238 91 240
rect 94 238 96 240
rect 99 238 101 240
rect 104 238 106 240
rect 109 238 111 240
rect 114 238 116 240
rect 183 238 185 240
rect 188 238 190 240
rect 193 238 195 240
rect 198 238 200 240
rect 203 238 205 240
rect 208 238 210 240
rect 213 238 215 240
rect 218 238 220 240
rect 223 238 225 240
rect 228 238 230 240
rect 233 238 235 240
rect 238 238 240 240
rect 243 238 245 240
rect 291 238 293 240
rect 296 238 298 240
rect 149 236 151 238
rect 271 235 273 237
rect 277 235 279 237
rect 3 233 5 235
rect 291 233 293 235
rect 296 233 298 235
rect 3 228 5 230
rect 18 229 20 231
rect 23 229 25 231
rect 55 230 57 232
rect 60 230 62 232
rect 70 230 72 232
rect 75 230 77 232
rect 85 230 87 232
rect 90 230 92 232
rect 100 230 102 232
rect 105 230 107 232
rect 115 230 117 232
rect 149 231 151 233
rect 183 230 185 232
rect 188 230 190 232
rect 198 230 200 232
rect 203 230 205 232
rect 213 230 215 232
rect 218 230 220 232
rect 228 230 230 232
rect 233 230 235 232
rect 243 230 245 232
rect 271 230 273 232
rect 277 230 279 232
rect 291 228 293 230
rect 296 228 298 230
rect 3 223 5 225
rect 55 224 57 226
rect 60 224 62 226
rect 70 224 72 226
rect 75 224 77 226
rect 85 224 87 226
rect 90 224 92 226
rect 100 224 102 226
rect 105 224 107 226
rect 115 224 117 226
rect 183 224 185 226
rect 188 224 190 226
rect 198 224 200 226
rect 203 224 205 226
rect 213 224 215 226
rect 218 224 220 226
rect 228 224 230 226
rect 233 224 235 226
rect 243 224 245 226
rect 277 225 279 227
rect 291 223 293 225
rect 296 223 298 225
rect 149 221 151 223
rect 3 218 5 220
rect 18 219 20 221
rect 23 219 25 221
rect 277 220 279 222
rect 291 218 293 220
rect 296 218 298 220
rect 149 216 151 218
rect 3 213 5 215
rect 18 214 20 216
rect 23 214 25 216
rect 33 214 35 216
rect 265 214 267 216
rect 277 215 279 217
rect 291 213 293 215
rect 296 213 298 215
rect 3 208 5 210
rect 18 209 20 211
rect 23 209 25 211
rect 33 209 35 211
rect 265 209 267 211
rect 277 210 279 212
rect 291 208 293 210
rect 296 208 298 210
rect 149 206 151 208
rect 3 203 5 205
rect 33 204 35 206
rect 265 204 267 206
rect 277 205 279 207
rect 291 203 293 205
rect 296 203 298 205
rect 149 201 151 203
rect 3 198 5 200
rect 18 199 20 201
rect 23 199 25 201
rect 33 199 35 201
rect 265 199 267 201
rect 277 200 279 202
rect 57 197 59 199
rect 62 197 64 199
rect 67 197 69 199
rect 72 197 74 199
rect 77 197 79 199
rect 82 197 84 199
rect 87 197 89 199
rect 92 197 94 199
rect 97 197 99 199
rect 102 197 104 199
rect 107 197 109 199
rect 112 197 114 199
rect 117 197 119 199
rect 181 197 183 199
rect 186 197 188 199
rect 191 197 193 199
rect 196 197 198 199
rect 201 197 203 199
rect 206 197 208 199
rect 211 197 213 199
rect 216 197 218 199
rect 221 197 223 199
rect 226 197 228 199
rect 231 197 233 199
rect 236 197 238 199
rect 241 197 243 199
rect 291 198 293 200
rect 296 198 298 200
rect 3 193 5 195
rect 18 194 20 196
rect 23 194 25 196
rect 33 194 35 196
rect 265 194 267 196
rect 277 195 279 197
rect 291 193 293 195
rect 296 193 298 195
rect 57 191 59 193
rect 62 191 64 193
rect 67 191 69 193
rect 72 191 74 193
rect 77 191 79 193
rect 82 191 84 193
rect 87 191 89 193
rect 92 191 94 193
rect 97 191 99 193
rect 102 191 104 193
rect 107 191 109 193
rect 112 191 114 193
rect 117 191 119 193
rect 149 191 151 193
rect 181 191 183 193
rect 186 191 188 193
rect 191 191 193 193
rect 196 191 198 193
rect 201 191 203 193
rect 206 191 208 193
rect 211 191 213 193
rect 216 191 218 193
rect 221 191 223 193
rect 226 191 228 193
rect 231 191 233 193
rect 236 191 238 193
rect 241 191 243 193
rect 3 188 5 190
rect 18 189 20 191
rect 23 189 25 191
rect 33 189 35 191
rect 265 189 267 191
rect 277 190 279 192
rect 291 188 293 190
rect 296 188 298 190
rect 149 186 151 188
rect 3 183 5 185
rect 33 184 35 186
rect 265 184 267 186
rect 277 185 279 187
rect 291 183 293 185
rect 296 183 298 185
rect 3 178 5 180
rect 18 179 20 181
rect 23 179 25 181
rect 33 179 35 181
rect 265 179 267 181
rect 277 180 279 182
rect 291 178 293 180
rect 296 178 298 180
rect 149 176 151 178
rect 3 173 5 175
rect 18 174 20 176
rect 23 174 25 176
rect 33 174 35 176
rect 265 174 267 176
rect 277 175 279 177
rect 291 173 293 175
rect 296 173 298 175
rect 149 171 151 173
rect 3 168 5 170
rect 18 169 20 171
rect 23 169 25 171
rect 33 169 35 171
rect 265 169 267 171
rect 277 170 279 172
rect 291 168 293 170
rect 296 168 298 170
rect 3 163 5 165
rect 33 164 35 166
rect 56 164 58 166
rect 61 164 63 166
rect 71 164 73 166
rect 76 164 78 166
rect 86 164 88 166
rect 91 164 93 166
rect 101 164 103 166
rect 106 164 108 166
rect 116 164 118 166
rect 182 164 184 166
rect 187 164 189 166
rect 197 164 199 166
rect 202 164 204 166
rect 212 164 214 166
rect 217 164 219 166
rect 227 164 229 166
rect 232 164 234 166
rect 242 164 244 166
rect 265 164 267 166
rect 277 165 279 167
rect 291 163 293 165
rect 296 163 298 165
rect 149 161 151 163
rect 3 158 5 160
rect 18 159 20 161
rect 23 159 25 161
rect 33 159 35 161
rect 56 158 58 160
rect 61 158 63 160
rect 71 158 73 160
rect 76 158 78 160
rect 86 158 88 160
rect 91 158 93 160
rect 101 158 103 160
rect 106 158 108 160
rect 116 158 118 160
rect 182 158 184 160
rect 187 158 189 160
rect 197 158 199 160
rect 202 158 204 160
rect 212 158 214 160
rect 217 158 219 160
rect 227 158 229 160
rect 232 158 234 160
rect 242 158 244 160
rect 265 159 267 161
rect 277 160 279 162
rect 291 158 293 160
rect 296 158 298 160
rect 149 156 151 158
rect 3 153 5 155
rect 18 154 20 156
rect 23 154 25 156
rect 33 154 35 156
rect 265 154 267 156
rect 277 155 279 157
rect 291 153 293 155
rect 296 153 298 155
rect 3 148 5 150
rect 18 149 20 151
rect 23 149 25 151
rect 33 149 35 151
rect 265 149 267 151
rect 277 150 279 152
rect 291 148 293 150
rect 296 148 298 150
rect 3 143 5 145
rect 33 144 35 146
rect 265 144 267 146
rect 277 145 279 147
rect 291 143 293 145
rect 296 143 298 145
rect 149 141 151 143
rect 3 138 5 140
rect 18 139 20 141
rect 23 139 25 141
rect 33 139 35 141
rect 265 139 267 141
rect 277 140 279 142
rect 291 138 293 140
rect 296 138 298 140
rect 3 133 5 135
rect 18 134 20 136
rect 23 134 25 136
rect 33 134 35 136
rect 265 134 267 136
rect 277 135 279 137
rect 291 133 293 135
rect 296 133 298 135
rect 57 131 59 133
rect 62 131 64 133
rect 67 131 69 133
rect 72 131 74 133
rect 77 131 79 133
rect 82 131 84 133
rect 87 131 89 133
rect 92 131 94 133
rect 97 131 99 133
rect 102 131 104 133
rect 107 131 109 133
rect 112 131 114 133
rect 117 131 119 133
rect 149 131 151 133
rect 181 131 183 133
rect 186 131 188 133
rect 191 131 193 133
rect 196 131 198 133
rect 201 131 203 133
rect 206 131 208 133
rect 211 131 213 133
rect 216 131 218 133
rect 221 131 223 133
rect 226 131 228 133
rect 231 131 233 133
rect 236 131 238 133
rect 241 131 243 133
rect 3 128 5 130
rect 18 129 20 131
rect 23 129 25 131
rect 33 129 35 131
rect 265 129 267 131
rect 277 130 279 132
rect 291 128 293 130
rect 296 128 298 130
rect 57 126 59 128
rect 62 126 64 128
rect 67 126 69 128
rect 72 126 74 128
rect 77 126 79 128
rect 82 126 84 128
rect 87 126 89 128
rect 92 126 94 128
rect 97 126 99 128
rect 102 126 104 128
rect 107 126 109 128
rect 112 126 114 128
rect 117 126 119 128
rect 149 126 151 128
rect 181 126 183 128
rect 186 126 188 128
rect 191 126 193 128
rect 196 126 198 128
rect 201 126 203 128
rect 206 126 208 128
rect 211 126 213 128
rect 216 126 218 128
rect 221 126 223 128
rect 226 126 228 128
rect 231 126 233 128
rect 236 126 238 128
rect 241 126 243 128
rect 3 123 5 125
rect 33 124 35 126
rect 265 124 267 126
rect 277 125 279 127
rect 291 123 293 125
rect 296 123 298 125
rect 3 118 5 120
rect 18 119 20 121
rect 23 119 25 121
rect 33 119 35 121
rect 265 119 267 121
rect 277 120 279 122
rect 291 118 293 120
rect 296 118 298 120
rect 149 116 151 118
rect 3 113 5 115
rect 18 114 20 116
rect 23 114 25 116
rect 33 114 35 116
rect 265 114 267 116
rect 277 115 279 117
rect 291 113 293 115
rect 296 113 298 115
rect 149 111 151 113
rect 3 108 5 110
rect 18 109 20 111
rect 23 109 25 111
rect 33 109 35 111
rect 265 109 267 111
rect 277 110 279 112
rect 291 108 293 110
rect 296 108 298 110
rect 3 103 5 105
rect 33 104 35 106
rect 265 104 267 106
rect 277 105 279 107
rect 291 103 293 105
rect 296 103 298 105
rect 149 101 151 103
rect 3 98 5 100
rect 18 99 20 101
rect 23 99 25 101
rect 33 99 35 101
rect 55 99 57 101
rect 60 99 62 101
rect 70 99 72 101
rect 75 99 77 101
rect 85 99 87 101
rect 90 99 92 101
rect 100 99 102 101
rect 105 99 107 101
rect 115 99 117 101
rect 183 99 185 101
rect 188 99 190 101
rect 198 99 200 101
rect 203 99 205 101
rect 213 99 215 101
rect 218 99 220 101
rect 228 99 230 101
rect 233 99 235 101
rect 243 99 245 101
rect 265 99 267 101
rect 277 100 279 102
rect 291 98 293 100
rect 296 98 298 100
rect 149 96 151 98
rect 3 93 5 95
rect 18 94 20 96
rect 23 94 25 96
rect 33 94 35 96
rect 55 93 57 95
rect 60 93 62 95
rect 70 93 72 95
rect 75 93 77 95
rect 85 93 87 95
rect 90 93 92 95
rect 100 93 102 95
rect 105 93 107 95
rect 115 93 117 95
rect 183 93 185 95
rect 188 93 190 95
rect 198 93 200 95
rect 203 93 205 95
rect 213 93 215 95
rect 218 93 220 95
rect 228 93 230 95
rect 233 93 235 95
rect 243 93 245 95
rect 265 94 267 96
rect 277 95 279 97
rect 291 93 293 95
rect 296 93 298 95
rect 3 88 5 90
rect 18 89 20 91
rect 23 89 25 91
rect 33 89 35 91
rect 265 89 267 91
rect 277 90 279 92
rect 291 88 293 90
rect 296 88 298 90
rect 149 86 151 88
rect 3 83 5 85
rect 33 84 35 86
rect 265 84 267 86
rect 277 85 279 87
rect 291 83 293 85
rect 296 83 298 85
rect 3 78 5 80
rect 18 79 20 81
rect 23 79 25 81
rect 33 79 35 81
rect 265 79 267 81
rect 277 80 279 82
rect 291 78 293 80
rect 296 78 298 80
rect 3 73 5 75
rect 18 74 20 76
rect 23 74 25 76
rect 33 74 35 76
rect 265 74 267 76
rect 277 75 279 77
rect 291 73 293 75
rect 296 73 298 75
rect 149 71 151 73
rect 3 68 5 70
rect 18 69 20 71
rect 23 69 25 71
rect 33 69 35 71
rect 265 69 267 71
rect 277 70 279 72
rect 291 68 293 70
rect 296 68 298 70
rect 57 66 59 68
rect 62 66 64 68
rect 67 66 69 68
rect 72 66 74 68
rect 77 66 79 68
rect 82 66 84 68
rect 87 66 89 68
rect 92 66 94 68
rect 97 66 99 68
rect 102 66 104 68
rect 107 66 109 68
rect 112 66 114 68
rect 117 66 119 68
rect 149 66 151 68
rect 181 66 183 68
rect 186 66 188 68
rect 191 66 193 68
rect 196 66 198 68
rect 201 66 203 68
rect 206 66 208 68
rect 211 66 213 68
rect 216 66 218 68
rect 221 66 223 68
rect 226 66 228 68
rect 231 66 233 68
rect 236 66 238 68
rect 241 66 243 68
rect 3 63 5 65
rect 33 64 35 66
rect 265 64 267 66
rect 277 65 279 67
rect 291 63 293 65
rect 296 63 298 65
rect 57 61 59 63
rect 62 61 64 63
rect 67 61 69 63
rect 72 61 74 63
rect 77 61 79 63
rect 82 61 84 63
rect 87 61 89 63
rect 92 61 94 63
rect 97 61 99 63
rect 102 61 104 63
rect 107 61 109 63
rect 112 61 114 63
rect 117 61 119 63
rect 181 61 183 63
rect 186 61 188 63
rect 191 61 193 63
rect 196 61 198 63
rect 201 61 203 63
rect 206 61 208 63
rect 211 61 213 63
rect 216 61 218 63
rect 221 61 223 63
rect 226 61 228 63
rect 231 61 233 63
rect 236 61 238 63
rect 241 61 243 63
rect 3 58 5 60
rect 18 59 20 61
rect 23 59 25 61
rect 33 59 35 61
rect 265 59 267 61
rect 277 60 279 62
rect 291 58 293 60
rect 296 58 298 60
rect 149 56 151 58
rect 3 53 5 55
rect 18 54 20 56
rect 23 54 25 56
rect 33 54 35 56
rect 265 54 267 56
rect 277 55 279 57
rect 291 53 293 55
rect 296 53 298 55
rect 3 48 5 50
rect 18 49 20 51
rect 23 49 25 51
rect 33 49 35 51
rect 265 49 267 51
rect 277 50 279 52
rect 291 48 293 50
rect 296 48 298 50
rect 3 43 5 45
rect 33 44 35 46
rect 265 44 267 46
rect 277 45 279 47
rect 291 43 293 45
rect 296 43 298 45
rect 3 38 5 40
rect 18 39 20 41
rect 23 39 25 41
rect 277 40 279 42
rect 291 38 293 40
rect 296 38 298 40
rect 3 33 5 35
rect 18 34 20 36
rect 23 34 25 36
rect 40 34 42 36
rect 54 34 56 36
rect 60 34 62 36
rect 65 34 67 36
rect 70 34 72 36
rect 75 34 77 36
rect 80 34 82 36
rect 85 34 87 36
rect 90 34 92 36
rect 95 34 97 36
rect 100 34 102 36
rect 105 34 107 36
rect 110 34 112 36
rect 115 34 117 36
rect 183 34 185 36
rect 188 34 190 36
rect 193 34 195 36
rect 198 34 200 36
rect 203 34 205 36
rect 208 34 210 36
rect 213 34 215 36
rect 218 34 220 36
rect 223 34 225 36
rect 228 34 230 36
rect 233 34 235 36
rect 238 34 240 36
rect 243 34 245 36
rect 277 35 279 37
rect 291 33 293 35
rect 296 33 298 35
rect 3 28 5 30
rect 40 28 42 30
rect 54 29 56 31
rect 277 30 279 32
rect 65 28 67 30
rect 75 28 77 30
rect 85 28 87 30
rect 95 28 97 30
rect 105 28 107 30
rect 115 28 117 30
rect 183 28 185 30
rect 193 28 195 30
rect 203 28 205 30
rect 213 28 215 30
rect 223 28 225 30
rect 233 28 235 30
rect 243 28 245 30
rect 18 26 20 28
rect 24 26 26 28
rect 29 26 31 28
rect 34 26 36 28
rect 264 27 266 29
rect 291 28 293 30
rect 296 28 298 30
rect 3 23 5 25
rect 54 24 56 26
rect 277 25 279 27
rect 65 23 67 25
rect 75 23 77 25
rect 85 23 87 25
rect 95 23 97 25
rect 105 23 107 25
rect 115 23 117 25
rect 183 23 185 25
rect 193 23 195 25
rect 203 23 205 25
rect 213 23 215 25
rect 223 23 225 25
rect 233 23 235 25
rect 243 23 245 25
rect 264 22 266 24
rect 291 23 293 25
rect 296 23 298 25
rect 3 18 5 20
rect 54 19 56 21
rect 277 20 279 22
rect 65 18 67 20
rect 75 18 77 20
rect 85 18 87 20
rect 95 18 97 20
rect 105 18 107 20
rect 115 18 117 20
rect 183 18 185 20
rect 193 18 195 20
rect 203 18 205 20
rect 213 18 215 20
rect 223 18 225 20
rect 233 18 235 20
rect 243 18 245 20
rect 24 16 26 18
rect 29 16 31 18
rect 34 16 36 18
rect 264 17 266 19
rect 291 18 293 20
rect 296 18 298 20
rect 277 15 279 17
rect 3 13 5 15
rect 291 13 293 15
rect 296 13 298 15
rect 3 8 5 10
rect 291 8 293 10
rect 296 8 298 10
rect 3 3 5 5
rect 9 3 11 5
rect 14 3 16 5
rect 19 3 21 5
rect 24 3 26 5
rect 29 3 31 5
rect 34 3 36 5
rect 39 3 41 5
rect 44 3 46 5
rect 49 3 51 5
rect 54 3 56 5
rect 59 3 61 5
rect 64 3 66 5
rect 69 3 71 5
rect 74 3 76 5
rect 79 3 81 5
rect 84 3 86 5
rect 89 3 91 5
rect 94 3 96 5
rect 99 3 101 5
rect 104 3 106 5
rect 109 3 111 5
rect 114 3 116 5
rect 119 3 121 5
rect 124 3 126 5
rect 129 3 131 5
rect 134 3 136 5
rect 139 3 141 5
rect 144 3 146 5
rect 149 3 151 5
rect 154 3 156 5
rect 159 3 161 5
rect 164 3 166 5
rect 169 3 171 5
rect 174 3 176 5
rect 179 3 181 5
rect 184 3 186 5
rect 189 3 191 5
rect 194 3 196 5
rect 199 3 201 5
rect 204 3 206 5
rect 209 3 211 5
rect 214 3 216 5
rect 219 3 221 5
rect 224 3 226 5
rect 229 3 231 5
rect 234 3 236 5
rect 239 3 241 5
rect 244 3 246 5
rect 249 3 251 5
rect 254 3 256 5
rect 259 3 261 5
rect 264 3 266 5
rect 269 3 271 5
rect 274 3 276 5
rect 279 3 281 5
rect 284 3 286 5
rect 291 3 293 5
rect 296 3 298 5
<< metal1 >>
rect 20 740 280 1000
rect 62 700 238 740
rect 102 690 198 700
rect 112 680 188 690
rect 0 658 116 669
rect 0 425 10 658
rect 14 617 117 655
rect 120 654 180 680
rect 184 658 300 669
rect 14 592 29 617
rect 32 595 36 614
rect 39 592 52 617
rect 120 612 143 654
rect 56 595 143 612
rect 14 552 117 592
rect 14 527 29 552
rect 32 530 36 549
rect 39 527 52 552
rect 120 548 143 595
rect 55 530 143 548
rect 14 488 117 527
rect 14 430 29 488
rect 32 436 36 481
rect 39 462 52 488
rect 120 483 143 530
rect 55 466 143 483
rect 39 439 116 462
rect 32 430 41 436
rect 44 430 116 439
rect 0 404 29 425
rect 0 354 11 404
rect 32 398 36 430
rect 39 410 115 425
rect 39 404 108 410
rect 120 407 143 466
rect 147 430 153 648
rect 157 612 180 654
rect 183 616 286 655
rect 157 595 244 612
rect 157 548 180 595
rect 248 590 261 616
rect 264 593 268 612
rect 271 590 286 616
rect 183 552 286 590
rect 157 530 244 548
rect 157 483 180 530
rect 248 527 261 552
rect 264 530 268 549
rect 271 527 286 552
rect 183 488 286 527
rect 157 466 244 483
rect 148 410 152 425
rect 157 407 180 466
rect 248 462 261 488
rect 184 439 261 462
rect 184 430 256 439
rect 264 436 268 484
rect 259 430 268 436
rect 271 430 286 488
rect 290 425 300 658
rect 184 410 300 425
rect 111 403 290 407
rect 32 393 41 398
rect 111 393 190 403
rect 37 390 41 393
rect 14 385 34 389
rect 37 387 131 390
rect 134 388 190 393
rect 193 390 208 400
rect 211 395 290 403
rect 211 390 228 395
rect 293 392 300 410
rect 127 385 131 387
rect 150 387 190 388
rect 211 387 215 390
rect 150 385 215 387
rect 14 360 18 385
rect 22 357 26 382
rect 19 354 26 357
rect 30 358 34 382
rect 39 381 123 384
rect 39 360 43 381
rect 30 354 35 358
rect 47 357 51 378
rect 0 341 6 354
rect 9 347 13 351
rect 19 348 22 354
rect 0 320 6 332
rect 9 327 12 347
rect 16 342 22 348
rect 25 347 29 351
rect 25 339 28 347
rect 32 339 35 354
rect 38 354 51 357
rect 55 355 59 381
rect 63 354 67 378
rect 71 355 75 381
rect 38 342 49 354
rect 64 352 67 354
rect 79 352 83 378
rect 87 355 91 381
rect 95 354 99 378
rect 103 356 107 381
rect 52 346 61 350
rect 20 335 29 339
rect 32 335 41 339
rect 9 323 13 327
rect 16 326 22 332
rect 19 320 22 326
rect 25 327 28 335
rect 25 323 29 327
rect 32 320 35 335
rect 0 272 11 320
rect 19 317 26 320
rect 14 273 18 314
rect 22 276 26 317
rect 30 316 35 320
rect 38 320 49 331
rect 53 327 56 346
rect 64 342 83 352
rect 86 347 95 351
rect 111 348 115 378
rect 119 360 123 381
rect 127 382 147 385
rect 158 383 215 385
rect 218 383 237 386
rect 127 357 131 382
rect 92 339 95 347
rect 98 342 115 348
rect 118 354 131 357
rect 135 357 139 379
rect 143 360 147 382
rect 151 357 155 382
rect 135 354 155 357
rect 80 335 89 339
rect 92 335 101 339
rect 52 323 61 327
rect 64 323 83 332
rect 86 327 89 335
rect 86 323 95 327
rect 98 326 115 332
rect 64 320 67 323
rect 38 317 51 320
rect 0 6 8 272
rect 14 270 27 273
rect 30 270 34 316
rect 39 273 43 314
rect 46 276 51 317
rect 55 274 59 320
rect 62 277 67 320
rect 55 273 60 274
rect 39 270 60 273
rect 63 272 67 277
rect 24 267 27 270
rect 57 269 60 270
rect 71 269 75 320
rect 78 272 83 323
rect 87 269 91 320
rect 94 272 99 318
rect 103 269 107 320
rect 111 276 115 326
rect 118 320 121 354
rect 151 353 155 354
rect 124 343 134 348
rect 137 347 146 351
rect 140 339 143 347
rect 124 335 133 339
rect 137 335 146 339
rect 127 327 130 335
rect 124 323 133 327
rect 136 326 148 332
rect 151 320 154 353
rect 118 317 139 320
rect 118 314 123 317
rect 119 273 123 314
rect 110 270 123 273
rect 127 275 131 313
rect 135 278 139 317
rect 143 317 154 320
rect 143 275 147 317
rect 127 271 147 275
rect 110 269 114 270
rect 11 263 20 267
rect 24 263 34 267
rect 45 263 54 267
rect 57 266 114 269
rect 127 267 131 271
rect 151 270 155 314
rect 117 264 131 267
rect 158 266 190 383
rect 218 380 221 383
rect 193 354 197 380
rect 201 377 221 380
rect 201 354 205 377
rect 194 348 197 354
rect 209 348 213 374
rect 194 336 213 348
rect 217 354 221 377
rect 224 354 229 380
rect 233 354 237 383
rect 249 383 285 386
rect 241 354 245 382
rect 249 354 253 383
rect 217 339 220 354
rect 224 347 227 354
rect 230 347 239 351
rect 242 348 245 354
rect 257 348 261 380
rect 223 343 227 347
rect 217 335 226 339
rect 194 326 213 332
rect 194 318 197 326
rect 11 13 14 263
rect 17 247 36 260
rect 17 221 36 243
rect 39 242 42 257
rect 39 232 43 242
rect 17 37 29 221
rect 39 217 42 232
rect 32 214 42 217
rect 32 43 36 214
rect 17 16 43 37
rect 23 14 40 16
rect 47 13 50 263
rect 57 260 114 263
rect 53 255 114 260
rect 53 253 108 255
rect 53 247 107 253
rect 117 251 120 264
rect 134 261 190 266
rect 111 247 120 251
rect 123 246 190 261
rect 193 260 197 318
rect 201 267 205 320
rect 209 272 213 326
rect 217 320 220 335
rect 223 327 227 331
rect 233 327 236 347
rect 242 342 261 348
rect 265 356 269 383
rect 224 320 227 327
rect 230 323 239 327
rect 242 326 261 332
rect 242 320 245 326
rect 217 267 221 320
rect 224 272 229 320
rect 233 267 237 320
rect 201 263 237 267
rect 193 247 230 260
rect 233 250 237 263
rect 241 260 245 320
rect 249 267 253 320
rect 257 272 261 326
rect 265 320 268 356
rect 272 355 277 380
rect 272 348 275 355
rect 281 354 285 383
rect 289 354 300 392
rect 271 342 275 348
rect 278 347 287 351
rect 280 339 283 347
rect 290 341 300 354
rect 277 335 286 339
rect 271 326 275 332
rect 280 327 283 335
rect 272 320 275 326
rect 278 323 287 327
rect 290 320 300 332
rect 265 267 269 320
rect 272 272 277 320
rect 281 267 285 320
rect 249 263 285 267
rect 240 253 254 260
rect 233 246 253 250
rect 123 244 176 246
rect 53 209 120 243
rect 123 205 143 244
rect 53 185 143 205
rect 53 143 120 182
rect 123 139 143 185
rect 56 120 143 139
rect 53 78 120 117
rect 123 74 143 120
rect 53 56 143 74
rect 53 18 119 52
rect 57 14 119 18
rect 123 49 143 56
rect 147 54 153 240
rect 157 205 176 244
rect 179 209 247 243
rect 157 185 247 205
rect 157 139 176 185
rect 180 143 247 182
rect 157 120 247 139
rect 157 74 176 120
rect 180 78 247 117
rect 157 56 247 74
rect 157 49 176 56
rect 11 9 20 13
rect 44 9 53 13
rect 123 12 176 49
rect 180 16 247 52
rect 180 14 241 16
rect 250 13 253 246
rect 244 9 253 13
rect 257 13 260 263
rect 289 260 300 320
rect 263 247 300 260
rect 263 232 267 242
rect 264 217 267 232
rect 270 229 286 243
rect 264 43 268 217
rect 271 37 286 229
rect 263 16 286 37
rect 269 14 286 16
rect 257 9 266 13
rect 289 8 300 247
rect 56 6 241 8
rect 269 6 300 8
rect 0 0 300 6
rect 111 -12 115 0
<< metal2 >>
rect 20 740 280 1000
rect 0 440 300 670
rect 0 439 29 440
rect 45 437 255 440
rect 271 439 300 440
rect 32 433 41 436
rect 259 433 268 436
rect 32 430 268 433
rect 36 429 268 430
rect 10 422 288 425
rect 0 368 300 422
rect 0 355 115 368
rect 119 360 139 364
rect 143 355 300 368
rect 0 343 300 355
rect 136 341 213 343
rect 242 342 261 343
rect 20 338 29 339
rect 92 338 101 339
rect 124 338 133 339
rect 20 335 133 338
rect 194 336 213 341
rect 217 338 226 339
rect 277 338 286 339
rect 217 335 286 338
rect 8 326 115 331
rect 136 329 213 332
rect 242 329 261 331
rect 136 326 261 329
rect 0 318 300 326
rect 0 306 131 318
rect 135 310 155 314
rect 159 306 300 318
rect 0 255 300 306
rect 0 253 108 255
rect 0 246 107 253
rect 111 242 120 251
rect 124 246 300 255
rect 39 238 267 242
rect 39 232 43 238
rect 0 228 35 230
rect 54 228 246 233
rect 263 232 267 238
rect 280 228 300 230
rect 0 23 300 228
rect 0 19 123 23
rect 0 0 7 19
rect 23 15 40 19
rect 11 -4 20 13
rect 24 0 40 15
rect 11 -6 29 -4
rect 14 -10 29 -6
rect 23 -19 29 -10
rect 44 -19 53 13
rect 57 0 123 19
rect 128 0 172 19
rect 176 17 300 23
rect 176 0 240 17
rect 263 16 267 17
rect 95 -12 99 0
rect 244 -19 253 13
rect 257 -19 266 13
rect 270 0 300 17
<< gv1 >>
rect 41 977 43 979
rect 53 977 55 979
rect 65 977 67 979
rect 77 977 79 979
rect 89 977 91 979
rect 101 977 103 979
rect 113 977 115 979
rect 125 977 127 979
rect 137 977 139 979
rect 149 977 151 979
rect 161 977 163 979
rect 173 977 175 979
rect 185 977 187 979
rect 197 977 199 979
rect 209 977 211 979
rect 221 977 223 979
rect 233 977 235 979
rect 245 977 247 979
rect 257 977 259 979
rect 41 965 43 967
rect 53 965 55 967
rect 65 965 67 967
rect 77 965 79 967
rect 89 965 91 967
rect 101 965 103 967
rect 113 965 115 967
rect 125 965 127 967
rect 137 965 139 967
rect 149 965 151 967
rect 161 965 163 967
rect 173 965 175 967
rect 185 965 187 967
rect 197 965 199 967
rect 209 965 211 967
rect 221 965 223 967
rect 233 965 235 967
rect 245 965 247 967
rect 257 965 259 967
rect 41 953 43 955
rect 53 953 55 955
rect 65 953 67 955
rect 77 953 79 955
rect 89 953 91 955
rect 101 953 103 955
rect 113 953 115 955
rect 125 953 127 955
rect 137 953 139 955
rect 149 953 151 955
rect 161 953 163 955
rect 173 953 175 955
rect 185 953 187 955
rect 197 953 199 955
rect 209 953 211 955
rect 221 953 223 955
rect 233 953 235 955
rect 245 953 247 955
rect 257 953 259 955
rect 41 941 43 943
rect 53 941 55 943
rect 65 941 67 943
rect 77 941 79 943
rect 89 941 91 943
rect 101 941 103 943
rect 113 941 115 943
rect 125 941 127 943
rect 137 941 139 943
rect 149 941 151 943
rect 161 941 163 943
rect 173 941 175 943
rect 185 941 187 943
rect 197 941 199 943
rect 209 941 211 943
rect 221 941 223 943
rect 233 941 235 943
rect 245 941 247 943
rect 257 941 259 943
rect 41 929 43 931
rect 53 929 55 931
rect 65 929 67 931
rect 77 929 79 931
rect 89 929 91 931
rect 101 929 103 931
rect 113 929 115 931
rect 125 929 127 931
rect 137 929 139 931
rect 149 929 151 931
rect 161 929 163 931
rect 173 929 175 931
rect 185 929 187 931
rect 197 929 199 931
rect 209 929 211 931
rect 221 929 223 931
rect 233 929 235 931
rect 245 929 247 931
rect 257 929 259 931
rect 41 917 43 919
rect 53 917 55 919
rect 65 917 67 919
rect 77 917 79 919
rect 89 917 91 919
rect 101 917 103 919
rect 113 917 115 919
rect 125 917 127 919
rect 137 917 139 919
rect 149 917 151 919
rect 161 917 163 919
rect 173 917 175 919
rect 185 917 187 919
rect 197 917 199 919
rect 209 917 211 919
rect 221 917 223 919
rect 233 917 235 919
rect 245 917 247 919
rect 257 917 259 919
rect 41 905 43 907
rect 53 905 55 907
rect 65 905 67 907
rect 77 905 79 907
rect 89 905 91 907
rect 101 905 103 907
rect 113 905 115 907
rect 125 905 127 907
rect 137 905 139 907
rect 149 905 151 907
rect 161 905 163 907
rect 173 905 175 907
rect 185 905 187 907
rect 197 905 199 907
rect 209 905 211 907
rect 221 905 223 907
rect 233 905 235 907
rect 245 905 247 907
rect 257 905 259 907
rect 41 893 43 895
rect 53 893 55 895
rect 65 893 67 895
rect 77 893 79 895
rect 89 893 91 895
rect 101 893 103 895
rect 113 893 115 895
rect 125 893 127 895
rect 137 893 139 895
rect 149 893 151 895
rect 161 893 163 895
rect 173 893 175 895
rect 185 893 187 895
rect 197 893 199 895
rect 209 893 211 895
rect 221 893 223 895
rect 233 893 235 895
rect 245 893 247 895
rect 257 893 259 895
rect 41 881 43 883
rect 53 881 55 883
rect 65 881 67 883
rect 77 881 79 883
rect 89 881 91 883
rect 101 881 103 883
rect 113 881 115 883
rect 125 881 127 883
rect 137 881 139 883
rect 149 881 151 883
rect 161 881 163 883
rect 173 881 175 883
rect 185 881 187 883
rect 197 881 199 883
rect 209 881 211 883
rect 221 881 223 883
rect 233 881 235 883
rect 245 881 247 883
rect 257 881 259 883
rect 41 869 43 871
rect 53 869 55 871
rect 65 869 67 871
rect 77 869 79 871
rect 89 869 91 871
rect 101 869 103 871
rect 113 869 115 871
rect 125 869 127 871
rect 137 869 139 871
rect 149 869 151 871
rect 161 869 163 871
rect 173 869 175 871
rect 185 869 187 871
rect 197 869 199 871
rect 209 869 211 871
rect 221 869 223 871
rect 233 869 235 871
rect 245 869 247 871
rect 257 869 259 871
rect 41 857 43 859
rect 53 857 55 859
rect 65 857 67 859
rect 77 857 79 859
rect 89 857 91 859
rect 101 857 103 859
rect 113 857 115 859
rect 125 857 127 859
rect 137 857 139 859
rect 149 857 151 859
rect 161 857 163 859
rect 173 857 175 859
rect 185 857 187 859
rect 197 857 199 859
rect 209 857 211 859
rect 221 857 223 859
rect 233 857 235 859
rect 245 857 247 859
rect 257 857 259 859
rect 41 845 43 847
rect 53 845 55 847
rect 65 845 67 847
rect 77 845 79 847
rect 89 845 91 847
rect 101 845 103 847
rect 113 845 115 847
rect 125 845 127 847
rect 137 845 139 847
rect 149 845 151 847
rect 161 845 163 847
rect 173 845 175 847
rect 185 845 187 847
rect 197 845 199 847
rect 209 845 211 847
rect 221 845 223 847
rect 233 845 235 847
rect 245 845 247 847
rect 257 845 259 847
rect 41 833 43 835
rect 53 833 55 835
rect 65 833 67 835
rect 77 833 79 835
rect 89 833 91 835
rect 101 833 103 835
rect 113 833 115 835
rect 125 833 127 835
rect 137 833 139 835
rect 149 833 151 835
rect 161 833 163 835
rect 173 833 175 835
rect 185 833 187 835
rect 197 833 199 835
rect 209 833 211 835
rect 221 833 223 835
rect 233 833 235 835
rect 245 833 247 835
rect 257 833 259 835
rect 41 821 43 823
rect 53 821 55 823
rect 65 821 67 823
rect 77 821 79 823
rect 89 821 91 823
rect 101 821 103 823
rect 113 821 115 823
rect 125 821 127 823
rect 137 821 139 823
rect 149 821 151 823
rect 161 821 163 823
rect 173 821 175 823
rect 185 821 187 823
rect 197 821 199 823
rect 209 821 211 823
rect 221 821 223 823
rect 233 821 235 823
rect 245 821 247 823
rect 257 821 259 823
rect 41 809 43 811
rect 53 809 55 811
rect 65 809 67 811
rect 77 809 79 811
rect 89 809 91 811
rect 101 809 103 811
rect 113 809 115 811
rect 125 809 127 811
rect 137 809 139 811
rect 149 809 151 811
rect 161 809 163 811
rect 173 809 175 811
rect 185 809 187 811
rect 197 809 199 811
rect 209 809 211 811
rect 221 809 223 811
rect 233 809 235 811
rect 245 809 247 811
rect 257 809 259 811
rect 41 797 43 799
rect 53 797 55 799
rect 65 797 67 799
rect 77 797 79 799
rect 89 797 91 799
rect 101 797 103 799
rect 113 797 115 799
rect 125 797 127 799
rect 137 797 139 799
rect 149 797 151 799
rect 161 797 163 799
rect 173 797 175 799
rect 185 797 187 799
rect 197 797 199 799
rect 209 797 211 799
rect 221 797 223 799
rect 233 797 235 799
rect 245 797 247 799
rect 257 797 259 799
rect 41 785 43 787
rect 53 785 55 787
rect 65 785 67 787
rect 77 785 79 787
rect 89 785 91 787
rect 101 785 103 787
rect 113 785 115 787
rect 125 785 127 787
rect 137 785 139 787
rect 149 785 151 787
rect 161 785 163 787
rect 173 785 175 787
rect 185 785 187 787
rect 197 785 199 787
rect 209 785 211 787
rect 221 785 223 787
rect 233 785 235 787
rect 245 785 247 787
rect 257 785 259 787
rect 41 773 43 775
rect 53 773 55 775
rect 65 773 67 775
rect 77 773 79 775
rect 89 773 91 775
rect 101 773 103 775
rect 113 773 115 775
rect 125 773 127 775
rect 137 773 139 775
rect 149 773 151 775
rect 161 773 163 775
rect 173 773 175 775
rect 185 773 187 775
rect 197 773 199 775
rect 209 773 211 775
rect 221 773 223 775
rect 233 773 235 775
rect 245 773 247 775
rect 257 773 259 775
rect 41 761 43 763
rect 53 761 55 763
rect 65 761 67 763
rect 77 761 79 763
rect 89 761 91 763
rect 101 761 103 763
rect 113 761 115 763
rect 125 761 127 763
rect 137 761 139 763
rect 149 761 151 763
rect 161 761 163 763
rect 173 761 175 763
rect 185 761 187 763
rect 197 761 199 763
rect 209 761 211 763
rect 221 761 223 763
rect 233 761 235 763
rect 245 761 247 763
rect 257 761 259 763
rect 15 651 17 653
rect 23 651 25 653
rect 28 651 30 653
rect 33 651 35 653
rect 38 651 40 653
rect 43 651 45 653
rect 48 651 50 653
rect 53 651 55 653
rect 58 651 60 653
rect 63 651 65 653
rect 68 651 70 653
rect 73 651 75 653
rect 78 651 80 653
rect 83 651 85 653
rect 88 651 90 653
rect 93 651 95 653
rect 98 651 100 653
rect 103 651 105 653
rect 108 651 110 653
rect 190 652 192 654
rect 195 652 197 654
rect 200 652 202 654
rect 205 652 207 654
rect 210 652 212 654
rect 215 652 217 654
rect 220 652 222 654
rect 225 652 227 654
rect 230 652 232 654
rect 235 652 237 654
rect 240 652 242 654
rect 245 652 247 654
rect 250 652 252 654
rect 255 652 257 654
rect 260 652 262 654
rect 265 652 267 654
rect 270 652 272 654
rect 275 652 277 654
rect 283 652 285 654
rect 15 646 17 648
rect 283 647 285 649
rect 15 641 17 643
rect 23 642 25 644
rect 31 642 33 644
rect 36 642 38 644
rect 41 642 43 644
rect 62 642 64 644
rect 77 642 79 644
rect 92 642 94 644
rect 107 642 109 644
rect 189 642 191 644
rect 204 642 206 644
rect 219 642 221 644
rect 234 642 236 644
rect 255 642 257 644
rect 260 642 262 644
rect 265 642 267 644
rect 272 642 274 644
rect 277 642 279 644
rect 283 642 285 644
rect 149 639 151 641
rect 15 636 17 638
rect 31 637 33 639
rect 36 637 38 639
rect 41 637 43 639
rect 62 637 64 639
rect 77 637 79 639
rect 92 637 94 639
rect 107 637 109 639
rect 189 637 191 639
rect 204 637 206 639
rect 219 637 221 639
rect 234 637 236 639
rect 255 637 257 639
rect 260 637 262 639
rect 265 637 267 639
rect 283 637 285 639
rect 15 631 17 633
rect 31 632 33 634
rect 36 632 38 634
rect 41 632 43 634
rect 62 632 64 634
rect 77 632 79 634
rect 92 632 94 634
rect 107 632 109 634
rect 189 632 191 634
rect 204 632 206 634
rect 219 632 221 634
rect 234 632 236 634
rect 255 632 257 634
rect 260 632 262 634
rect 265 632 267 634
rect 283 632 285 634
rect 15 626 17 628
rect 283 627 285 629
rect 15 621 17 623
rect 21 622 23 624
rect 26 622 28 624
rect 33 622 35 624
rect 265 622 267 624
rect 272 622 274 624
rect 277 622 279 624
rect 283 622 285 624
rect 42 618 44 620
rect 47 618 49 620
rect 53 619 55 621
rect 58 619 60 621
rect 63 619 65 621
rect 68 619 70 621
rect 73 619 75 621
rect 78 619 80 621
rect 83 619 85 621
rect 88 619 90 621
rect 93 619 95 621
rect 98 619 100 621
rect 103 619 105 621
rect 108 619 110 621
rect 113 619 115 621
rect 149 619 151 621
rect 187 619 189 621
rect 192 619 194 621
rect 197 619 199 621
rect 202 619 204 621
rect 207 619 209 621
rect 212 619 214 621
rect 217 619 219 621
rect 222 619 224 621
rect 227 619 229 621
rect 232 619 234 621
rect 237 619 239 621
rect 242 619 244 621
rect 15 616 17 618
rect 250 617 252 619
rect 255 617 257 619
rect 283 617 285 619
rect 42 613 44 615
rect 47 613 49 615
rect 15 611 17 613
rect 250 612 252 614
rect 255 612 257 614
rect 283 612 285 614
rect 42 608 44 610
rect 47 608 49 610
rect 15 606 17 608
rect 250 607 252 609
rect 255 607 257 609
rect 283 607 285 609
rect 15 601 17 603
rect 21 602 23 604
rect 26 602 28 604
rect 42 603 44 605
rect 47 603 49 605
rect 250 602 252 604
rect 255 602 257 604
rect 272 602 274 604
rect 277 602 279 604
rect 283 602 285 604
rect 42 598 44 600
rect 47 598 49 600
rect 149 599 151 601
rect 15 596 17 598
rect 250 597 252 599
rect 255 597 257 599
rect 283 597 285 599
rect 42 593 44 595
rect 47 593 49 595
rect 15 591 17 593
rect 250 592 252 594
rect 255 592 257 594
rect 283 592 285 594
rect 42 588 44 590
rect 47 588 49 590
rect 15 586 17 588
rect 33 586 35 588
rect 53 587 55 589
rect 58 587 60 589
rect 63 587 65 589
rect 68 587 70 589
rect 73 587 75 589
rect 78 587 80 589
rect 83 587 85 589
rect 88 587 90 589
rect 93 587 95 589
rect 98 587 100 589
rect 103 587 105 589
rect 108 587 110 589
rect 113 587 115 589
rect 187 586 189 588
rect 192 586 194 588
rect 197 586 199 588
rect 202 586 204 588
rect 207 586 209 588
rect 212 586 214 588
rect 217 586 219 588
rect 222 586 224 588
rect 227 586 229 588
rect 232 586 234 588
rect 237 586 239 588
rect 242 586 244 588
rect 250 587 252 589
rect 255 587 257 589
rect 283 587 285 589
rect 265 585 267 587
rect 15 581 17 583
rect 21 582 23 584
rect 26 582 28 584
rect 33 581 35 583
rect 272 582 274 584
rect 277 582 279 584
rect 283 582 285 584
rect 149 579 151 581
rect 265 580 267 582
rect 15 576 17 578
rect 33 576 35 578
rect 283 577 285 579
rect 265 575 267 577
rect 42 573 44 575
rect 47 573 49 575
rect 52 573 54 575
rect 57 573 59 575
rect 72 573 74 575
rect 87 573 89 575
rect 102 573 104 575
rect 195 573 197 575
rect 210 573 212 575
rect 225 573 227 575
rect 240 573 242 575
rect 245 573 247 575
rect 250 573 252 575
rect 255 573 257 575
rect 15 571 17 573
rect 33 571 35 573
rect 283 572 285 574
rect 265 570 267 572
rect 15 566 17 568
rect 33 566 35 568
rect 42 567 44 569
rect 47 567 49 569
rect 52 567 54 569
rect 57 567 59 569
rect 72 567 74 569
rect 87 567 89 569
rect 102 567 104 569
rect 195 567 197 569
rect 210 567 212 569
rect 225 567 227 569
rect 240 567 242 569
rect 245 567 247 569
rect 250 567 252 569
rect 255 567 257 569
rect 283 567 285 569
rect 265 565 267 567
rect 15 561 17 563
rect 21 562 23 564
rect 26 562 28 564
rect 33 561 35 563
rect 272 562 274 564
rect 277 562 279 564
rect 283 562 285 564
rect 149 559 151 561
rect 265 560 267 562
rect 15 556 17 558
rect 33 556 35 558
rect 283 557 285 559
rect 43 553 45 555
rect 48 553 50 555
rect 56 553 58 555
rect 61 553 63 555
rect 66 553 68 555
rect 71 553 73 555
rect 76 553 78 555
rect 81 553 83 555
rect 86 553 88 555
rect 91 553 93 555
rect 96 553 98 555
rect 101 553 103 555
rect 106 553 108 555
rect 111 553 113 555
rect 187 554 189 556
rect 192 554 194 556
rect 197 554 199 556
rect 202 554 204 556
rect 207 554 209 556
rect 212 554 214 556
rect 217 554 219 556
rect 222 554 224 556
rect 227 554 229 556
rect 232 554 234 556
rect 237 554 239 556
rect 242 554 244 556
rect 265 555 267 557
rect 250 553 252 555
rect 255 553 257 555
rect 15 551 17 553
rect 283 552 285 554
rect 43 548 45 550
rect 48 548 50 550
rect 250 548 252 550
rect 255 548 257 550
rect 15 546 17 548
rect 283 547 285 549
rect 15 541 17 543
rect 21 542 23 544
rect 26 542 28 544
rect 43 543 45 545
rect 48 543 50 545
rect 250 543 252 545
rect 255 543 257 545
rect 272 542 274 544
rect 277 542 279 544
rect 283 542 285 544
rect 43 538 45 540
rect 48 538 50 540
rect 149 539 151 541
rect 250 538 252 540
rect 255 538 257 540
rect 15 536 17 538
rect 283 537 285 539
rect 43 533 45 535
rect 48 533 50 535
rect 250 533 252 535
rect 255 533 257 535
rect 15 531 17 533
rect 283 532 285 534
rect 43 528 45 530
rect 48 528 50 530
rect 250 528 252 530
rect 255 528 257 530
rect 15 526 17 528
rect 283 527 285 529
rect 15 521 17 523
rect 21 522 23 524
rect 26 522 28 524
rect 43 523 45 525
rect 48 523 50 525
rect 56 523 58 525
rect 61 523 63 525
rect 66 523 68 525
rect 71 523 73 525
rect 76 523 78 525
rect 81 523 83 525
rect 86 523 88 525
rect 91 523 93 525
rect 96 523 98 525
rect 101 523 103 525
rect 106 523 108 525
rect 111 523 113 525
rect 187 523 189 525
rect 192 523 194 525
rect 197 523 199 525
rect 202 523 204 525
rect 207 523 209 525
rect 212 523 214 525
rect 217 523 219 525
rect 222 523 224 525
rect 227 523 229 525
rect 232 523 234 525
rect 237 523 239 525
rect 242 523 244 525
rect 250 523 252 525
rect 255 523 257 525
rect 33 521 35 523
rect 265 521 267 523
rect 272 522 274 524
rect 277 522 279 524
rect 283 522 285 524
rect 149 519 151 521
rect 15 516 17 518
rect 33 516 35 518
rect 265 516 267 518
rect 283 517 285 519
rect 15 511 17 513
rect 33 511 35 513
rect 265 511 267 513
rect 283 512 285 514
rect 42 509 44 511
rect 47 509 49 511
rect 52 509 54 511
rect 57 509 59 511
rect 72 509 74 511
rect 87 509 89 511
rect 102 509 104 511
rect 194 509 196 511
rect 209 509 211 511
rect 224 509 226 511
rect 239 509 241 511
rect 244 509 246 511
rect 249 509 251 511
rect 254 509 256 511
rect 15 506 17 508
rect 33 506 35 508
rect 265 506 267 508
rect 283 507 285 509
rect 15 501 17 503
rect 21 502 23 504
rect 26 502 28 504
rect 42 503 44 505
rect 47 503 49 505
rect 52 503 54 505
rect 57 503 59 505
rect 72 503 74 505
rect 87 503 89 505
rect 102 503 104 505
rect 194 503 196 505
rect 209 503 211 505
rect 224 503 226 505
rect 239 503 241 505
rect 244 503 246 505
rect 249 503 251 505
rect 254 503 256 505
rect 33 501 35 503
rect 265 501 267 503
rect 272 502 274 504
rect 277 502 279 504
rect 283 502 285 504
rect 149 499 151 501
rect 15 496 17 498
rect 33 496 35 498
rect 265 496 267 498
rect 283 497 285 499
rect 15 491 17 493
rect 33 491 35 493
rect 43 489 45 491
rect 48 489 50 491
rect 56 490 58 492
rect 61 490 63 492
rect 66 490 68 492
rect 71 490 73 492
rect 76 490 78 492
rect 81 490 83 492
rect 86 490 88 492
rect 91 490 93 492
rect 96 490 98 492
rect 101 490 103 492
rect 106 490 108 492
rect 111 490 113 492
rect 185 490 187 492
rect 190 490 192 492
rect 195 490 197 492
rect 200 490 202 492
rect 205 490 207 492
rect 210 490 212 492
rect 215 490 217 492
rect 220 490 222 492
rect 225 490 227 492
rect 230 490 232 492
rect 235 490 237 492
rect 240 490 242 492
rect 245 490 247 492
rect 265 491 267 493
rect 283 492 285 494
rect 251 489 253 491
rect 256 489 258 491
rect 15 486 17 488
rect 283 487 285 489
rect 43 484 45 486
rect 48 484 50 486
rect 251 484 253 486
rect 256 484 258 486
rect 15 481 17 483
rect 21 482 23 484
rect 26 482 28 484
rect 272 482 274 484
rect 277 482 279 484
rect 283 482 285 484
rect 43 479 45 481
rect 48 479 50 481
rect 149 479 151 481
rect 251 479 253 481
rect 256 479 258 481
rect 15 476 17 478
rect 283 477 285 479
rect 43 474 45 476
rect 48 474 50 476
rect 251 474 253 476
rect 256 474 258 476
rect 15 471 17 473
rect 283 472 285 474
rect 43 469 45 471
rect 48 469 50 471
rect 251 469 253 471
rect 256 469 258 471
rect 15 466 17 468
rect 283 467 285 469
rect 43 464 45 466
rect 48 464 50 466
rect 251 464 253 466
rect 256 464 258 466
rect 15 461 17 463
rect 21 462 23 464
rect 26 462 28 464
rect 272 462 274 464
rect 277 462 279 464
rect 283 462 285 464
rect 43 459 45 461
rect 48 459 50 461
rect 55 458 57 460
rect 60 458 62 460
rect 65 458 67 460
rect 70 458 72 460
rect 75 458 77 460
rect 80 458 82 460
rect 85 458 87 460
rect 90 458 92 460
rect 95 458 97 460
rect 100 458 102 460
rect 105 458 107 460
rect 110 458 112 460
rect 149 459 151 461
rect 188 458 190 460
rect 193 458 195 460
rect 198 458 200 460
rect 203 458 205 460
rect 208 458 210 460
rect 213 458 215 460
rect 218 458 220 460
rect 223 458 225 460
rect 228 458 230 460
rect 233 458 235 460
rect 238 458 240 460
rect 243 458 245 460
rect 251 459 253 461
rect 256 459 258 461
rect 15 456 17 458
rect 283 457 285 459
rect 15 451 17 453
rect 283 452 285 454
rect 15 446 17 448
rect 283 447 285 449
rect 41 444 43 446
rect 46 444 48 446
rect 52 444 54 446
rect 57 444 59 446
rect 72 444 74 446
rect 87 444 89 446
rect 102 444 104 446
rect 195 444 197 446
rect 210 444 212 446
rect 225 444 227 446
rect 240 444 242 446
rect 246 444 248 446
rect 251 444 253 446
rect 257 444 259 446
rect 15 441 17 443
rect 21 442 23 444
rect 26 442 28 444
rect 272 442 274 444
rect 277 442 279 444
rect 283 442 285 444
rect 47 438 49 440
rect 57 438 59 440
rect 72 438 74 440
rect 87 438 89 440
rect 102 438 104 440
rect 149 439 151 441
rect 195 438 197 440
rect 210 438 212 440
rect 225 438 227 440
rect 240 438 242 440
rect 250 438 252 440
rect 33 432 35 434
rect 38 432 40 434
rect 260 432 262 434
rect 265 432 267 434
rect 16 422 18 424
rect 21 422 23 424
rect 26 422 28 424
rect 40 422 42 424
rect 45 422 47 424
rect 50 422 52 424
rect 55 422 57 424
rect 60 422 62 424
rect 65 422 67 424
rect 70 422 72 424
rect 75 422 77 424
rect 80 422 82 424
rect 85 422 87 424
rect 90 422 92 424
rect 95 422 97 424
rect 100 422 102 424
rect 105 422 107 424
rect 110 422 112 424
rect 149 422 151 424
rect 185 422 187 424
rect 190 422 192 424
rect 195 422 197 424
rect 200 422 202 424
rect 205 422 207 424
rect 210 422 212 424
rect 215 422 217 424
rect 220 422 222 424
rect 225 422 227 424
rect 230 422 232 424
rect 235 422 237 424
rect 240 422 242 424
rect 245 422 247 424
rect 250 422 252 424
rect 255 422 257 424
rect 260 422 262 424
rect 265 422 267 424
rect 270 422 272 424
rect 275 422 277 424
rect 280 422 282 424
rect 285 422 287 424
rect 296 408 298 410
rect 8 406 10 408
rect 14 406 16 408
rect 19 406 21 408
rect 24 406 26 408
rect 40 406 42 408
rect 45 406 47 408
rect 50 406 52 408
rect 55 406 57 408
rect 60 406 62 408
rect 65 406 67 408
rect 70 406 72 408
rect 75 406 77 408
rect 80 406 82 408
rect 85 406 87 408
rect 90 406 92 408
rect 95 406 97 408
rect 100 406 102 408
rect 105 406 107 408
rect 8 401 10 403
rect 296 398 298 400
rect 8 396 10 398
rect 8 390 10 392
rect 290 389 292 391
rect 296 388 298 390
rect 8 385 10 387
rect 8 380 10 382
rect 296 378 298 380
rect 8 375 10 377
rect 23 372 25 374
rect 194 372 196 374
rect 226 372 228 374
rect 242 372 244 374
rect 258 372 260 374
rect 274 372 276 374
rect 290 372 292 374
rect 8 370 10 372
rect 48 370 50 372
rect 64 370 66 372
rect 80 370 82 372
rect 96 370 98 372
rect 112 370 114 372
rect 296 368 298 370
rect 8 365 10 367
rect 23 362 25 364
rect 8 360 10 362
rect 48 360 50 362
rect 64 360 66 362
rect 80 360 82 362
rect 96 360 98 362
rect 112 360 114 362
rect 120 361 122 363
rect 136 361 138 363
rect 194 362 196 364
rect 210 361 212 363
rect 226 362 228 364
rect 242 362 244 364
rect 258 362 260 364
rect 274 362 276 364
rect 290 362 292 364
rect 296 358 298 360
rect 8 355 10 357
rect 291 348 293 350
rect 296 348 298 350
rect 104 344 106 346
rect 131 344 133 346
rect 253 343 255 345
rect 21 336 23 338
rect 26 336 28 338
rect 93 336 95 338
rect 98 336 100 338
rect 125 336 127 338
rect 130 336 132 338
rect 195 337 197 339
rect 200 337 202 339
rect 205 337 207 339
rect 210 337 212 339
rect 218 336 220 338
rect 223 336 225 338
rect 278 336 280 338
rect 283 336 285 338
rect 70 328 72 330
rect 105 328 107 330
rect 143 328 145 330
rect 205 328 207 330
rect 253 328 255 330
rect 80 318 82 320
rect 296 318 298 320
rect 8 315 10 317
rect 23 312 25 314
rect 48 312 50 314
rect 112 312 114 314
rect 296 313 298 315
rect 8 310 10 312
rect 136 311 138 313
rect 152 311 154 313
rect 64 308 66 310
rect 80 308 82 310
rect 96 308 98 310
rect 194 308 196 310
rect 210 308 212 310
rect 226 308 228 310
rect 242 308 244 310
rect 258 308 260 310
rect 274 308 276 310
rect 296 308 298 310
rect 8 305 10 307
rect 23 302 25 304
rect 48 302 50 304
rect 112 302 114 304
rect 296 303 298 305
rect 8 300 10 302
rect 64 298 66 300
rect 80 298 82 300
rect 96 298 98 300
rect 194 298 196 300
rect 210 298 212 300
rect 226 298 228 300
rect 242 298 244 300
rect 258 298 260 300
rect 274 298 276 300
rect 296 298 298 300
rect 8 295 10 297
rect 23 292 25 294
rect 48 292 50 294
rect 112 292 114 294
rect 194 293 196 295
rect 210 293 212 295
rect 226 293 228 295
rect 242 293 244 295
rect 258 293 260 295
rect 274 293 276 295
rect 296 293 298 295
rect 8 290 10 292
rect 64 288 66 290
rect 80 288 82 290
rect 96 288 98 290
rect 296 288 298 290
rect 8 285 10 287
rect 23 282 25 284
rect 48 282 50 284
rect 112 282 114 284
rect 296 283 298 285
rect 8 280 10 282
rect 64 278 66 280
rect 80 278 82 280
rect 96 278 98 280
rect 194 278 196 280
rect 210 278 212 280
rect 226 278 228 280
rect 242 278 244 280
rect 258 278 260 280
rect 274 278 276 280
rect 296 278 298 280
rect 8 275 10 277
rect 296 273 298 275
rect 296 268 298 270
rect 296 263 298 265
rect 296 258 298 260
rect 18 248 20 250
rect 23 248 25 250
rect 28 248 30 250
rect 33 248 35 250
rect 54 248 56 250
rect 59 248 61 250
rect 64 248 66 250
rect 69 248 71 250
rect 74 248 76 250
rect 79 248 81 250
rect 84 248 86 250
rect 89 248 91 250
rect 94 248 96 250
rect 99 248 101 250
rect 104 248 106 250
rect 112 248 114 250
rect 117 248 119 250
rect 195 248 197 250
rect 200 248 202 250
rect 205 248 207 250
rect 210 248 212 250
rect 215 248 217 250
rect 220 248 222 250
rect 225 248 227 250
rect 264 248 266 250
rect 269 248 271 250
rect 274 248 276 250
rect 279 248 281 250
rect 284 248 286 250
rect 40 239 42 241
rect 264 239 266 241
rect 40 233 42 235
rect 264 233 266 235
rect 65 230 67 232
rect 80 230 82 232
rect 95 230 97 232
rect 110 230 112 232
rect 193 230 195 232
rect 208 230 210 232
rect 223 230 225 232
rect 238 230 240 232
rect 149 226 151 228
rect 18 224 20 226
rect 23 224 25 226
rect 33 223 35 225
rect 65 224 67 226
rect 80 224 82 226
rect 95 224 97 226
rect 110 224 112 226
rect 193 224 195 226
rect 208 224 210 226
rect 223 224 225 226
rect 238 224 240 226
rect 272 225 274 227
rect 283 225 285 227
rect 272 220 274 222
rect 283 220 285 222
rect 272 215 274 217
rect 283 215 285 217
rect 55 211 57 213
rect 60 211 62 213
rect 65 211 67 213
rect 70 211 72 213
rect 75 211 77 213
rect 80 211 82 213
rect 85 211 87 213
rect 90 211 92 213
rect 95 211 97 213
rect 100 211 102 213
rect 105 211 107 213
rect 110 211 112 213
rect 115 211 117 213
rect 149 211 151 213
rect 183 211 185 213
rect 188 211 190 213
rect 193 211 195 213
rect 198 211 200 213
rect 203 211 205 213
rect 208 211 210 213
rect 213 211 215 213
rect 218 211 220 213
rect 223 211 225 213
rect 228 211 230 213
rect 233 211 235 213
rect 238 211 240 213
rect 243 211 245 213
rect 272 210 274 212
rect 283 210 285 212
rect 18 204 20 206
rect 23 204 25 206
rect 272 205 274 207
rect 283 205 285 207
rect 272 200 274 202
rect 283 200 285 202
rect 149 196 151 198
rect 272 195 274 197
rect 283 195 285 197
rect 272 190 274 192
rect 283 190 285 192
rect 18 184 20 186
rect 23 184 25 186
rect 272 185 274 187
rect 283 185 285 187
rect 149 181 151 183
rect 272 180 274 182
rect 283 180 285 182
rect 57 178 59 180
rect 62 178 64 180
rect 67 178 69 180
rect 72 178 74 180
rect 77 178 79 180
rect 82 178 84 180
rect 87 178 89 180
rect 92 178 94 180
rect 97 178 99 180
rect 102 178 104 180
rect 107 178 109 180
rect 112 178 114 180
rect 117 178 119 180
rect 183 178 185 180
rect 188 178 190 180
rect 193 178 195 180
rect 198 178 200 180
rect 203 178 205 180
rect 208 178 210 180
rect 213 178 215 180
rect 218 178 220 180
rect 223 178 225 180
rect 228 178 230 180
rect 233 178 235 180
rect 238 178 240 180
rect 243 178 245 180
rect 272 175 274 177
rect 283 175 285 177
rect 272 170 274 172
rect 283 170 285 172
rect 149 166 151 168
rect 18 164 20 166
rect 23 164 25 166
rect 66 164 68 166
rect 81 164 83 166
rect 96 164 98 166
rect 111 164 113 166
rect 192 164 194 166
rect 207 164 209 166
rect 222 164 224 166
rect 237 164 239 166
rect 272 165 274 167
rect 283 165 285 167
rect 272 160 274 162
rect 283 160 285 162
rect 66 158 68 160
rect 81 158 83 160
rect 96 158 98 160
rect 111 158 113 160
rect 192 158 194 160
rect 207 158 209 160
rect 222 158 224 160
rect 237 158 239 160
rect 272 155 274 157
rect 283 155 285 157
rect 149 151 151 153
rect 272 150 274 152
rect 283 150 285 152
rect 18 144 20 146
rect 23 144 25 146
rect 56 145 58 147
rect 61 145 63 147
rect 66 145 68 147
rect 71 145 73 147
rect 76 145 78 147
rect 81 145 83 147
rect 86 145 88 147
rect 91 145 93 147
rect 96 145 98 147
rect 101 145 103 147
rect 106 145 108 147
rect 111 145 113 147
rect 116 145 118 147
rect 182 145 184 147
rect 187 145 189 147
rect 192 145 194 147
rect 197 145 199 147
rect 202 145 204 147
rect 207 145 209 147
rect 212 145 214 147
rect 217 145 219 147
rect 222 145 224 147
rect 227 145 229 147
rect 232 145 234 147
rect 237 145 239 147
rect 242 145 244 147
rect 272 145 274 147
rect 283 145 285 147
rect 272 140 274 142
rect 283 140 285 142
rect 149 136 151 138
rect 272 135 274 137
rect 283 135 285 137
rect 272 130 274 132
rect 283 130 285 132
rect 18 124 20 126
rect 23 124 25 126
rect 272 125 274 127
rect 283 125 285 127
rect 149 121 151 123
rect 272 120 274 122
rect 283 120 285 122
rect 272 115 274 117
rect 283 115 285 117
rect 56 113 58 115
rect 61 113 63 115
rect 66 113 68 115
rect 71 113 73 115
rect 76 113 78 115
rect 81 113 83 115
rect 86 113 88 115
rect 91 113 93 115
rect 96 113 98 115
rect 101 113 103 115
rect 106 113 108 115
rect 111 113 113 115
rect 116 113 118 115
rect 183 112 185 114
rect 188 112 190 114
rect 193 112 195 114
rect 198 112 200 114
rect 203 112 205 114
rect 208 112 210 114
rect 213 112 215 114
rect 218 112 220 114
rect 223 112 225 114
rect 228 112 230 114
rect 233 112 235 114
rect 238 112 240 114
rect 243 112 245 114
rect 272 110 274 112
rect 283 110 285 112
rect 149 106 151 108
rect 18 104 20 106
rect 23 104 25 106
rect 272 105 274 107
rect 283 105 285 107
rect 65 99 67 101
rect 80 99 82 101
rect 95 99 97 101
rect 110 99 112 101
rect 193 99 195 101
rect 208 99 210 101
rect 223 99 225 101
rect 238 99 240 101
rect 272 100 274 102
rect 283 100 285 102
rect 272 95 274 97
rect 283 95 285 97
rect 65 93 67 95
rect 80 93 82 95
rect 95 93 97 95
rect 110 93 112 95
rect 193 93 195 95
rect 208 93 210 95
rect 223 93 225 95
rect 238 93 240 95
rect 149 91 151 93
rect 272 90 274 92
rect 283 90 285 92
rect 18 84 20 86
rect 23 84 25 86
rect 272 85 274 87
rect 283 85 285 87
rect 56 81 58 83
rect 61 81 63 83
rect 66 81 68 83
rect 71 81 73 83
rect 76 81 78 83
rect 81 81 83 83
rect 86 81 88 83
rect 91 81 93 83
rect 96 81 98 83
rect 101 81 103 83
rect 106 81 108 83
rect 111 81 113 83
rect 116 81 118 83
rect 183 81 185 83
rect 188 81 190 83
rect 193 81 195 83
rect 198 81 200 83
rect 203 81 205 83
rect 208 81 210 83
rect 213 81 215 83
rect 218 81 220 83
rect 223 81 225 83
rect 228 81 230 83
rect 233 81 235 83
rect 238 81 240 83
rect 243 81 245 83
rect 272 80 274 82
rect 283 80 285 82
rect 149 76 151 78
rect 272 75 274 77
rect 283 75 285 77
rect 272 70 274 72
rect 283 70 285 72
rect 18 64 20 66
rect 23 64 25 66
rect 272 65 274 67
rect 283 65 285 67
rect 149 61 151 63
rect 272 60 274 62
rect 283 60 285 62
rect 272 55 274 57
rect 283 55 285 57
rect 272 50 274 52
rect 283 50 285 52
rect 55 48 57 50
rect 60 48 62 50
rect 65 48 67 50
rect 70 48 72 50
rect 75 48 77 50
rect 80 48 82 50
rect 85 48 87 50
rect 90 48 92 50
rect 95 48 97 50
rect 100 48 102 50
rect 105 48 107 50
rect 110 48 112 50
rect 115 48 117 50
rect 183 48 185 50
rect 188 48 190 50
rect 193 48 195 50
rect 198 48 200 50
rect 203 48 205 50
rect 208 48 210 50
rect 213 48 215 50
rect 218 48 220 50
rect 223 48 225 50
rect 228 48 230 50
rect 233 48 235 50
rect 238 48 240 50
rect 243 48 245 50
rect 18 44 20 46
rect 23 44 25 46
rect 272 45 274 47
rect 283 45 285 47
rect 272 40 274 42
rect 283 40 285 42
rect 272 35 274 37
rect 283 35 285 37
rect 33 33 35 35
rect 265 33 267 35
rect 272 30 274 32
rect 283 30 285 32
rect 60 28 62 30
rect 70 28 72 30
rect 80 28 82 30
rect 90 28 92 30
rect 100 28 102 30
rect 110 28 112 30
rect 188 28 190 30
rect 198 28 200 30
rect 208 28 210 30
rect 218 28 220 30
rect 228 28 230 30
rect 238 28 240 30
rect 40 24 42 26
rect 272 25 274 27
rect 283 25 285 27
rect 60 23 62 25
rect 70 23 72 25
rect 80 23 82 25
rect 90 23 92 25
rect 100 23 102 25
rect 110 23 112 25
rect 188 23 190 25
rect 198 23 200 25
rect 208 23 210 25
rect 218 23 220 25
rect 228 23 230 25
rect 238 23 240 25
rect 18 21 20 23
rect 24 21 26 23
rect 29 21 31 23
rect 34 21 36 23
rect 272 20 274 22
rect 283 20 285 22
rect 60 18 62 20
rect 70 18 72 20
rect 80 18 82 20
rect 90 18 92 20
rect 100 18 102 20
rect 110 18 112 20
rect 188 18 190 20
rect 198 18 200 20
rect 208 18 210 20
rect 218 18 220 20
rect 228 18 230 20
rect 238 18 240 20
rect 129 16 131 18
rect 134 16 136 18
rect 139 16 141 18
rect 144 16 146 18
rect 149 16 151 18
rect 154 16 156 18
rect 159 16 161 18
rect 164 16 166 18
rect 169 16 171 18
rect 272 15 274 17
rect 283 15 285 17
rect 12 10 14 12
rect 17 10 19 12
rect 45 10 47 12
rect 50 10 52 12
rect 245 10 247 12
rect 250 10 252 12
rect 258 10 260 12
rect 263 10 265 12
<< metal3 >>
rect 23 743 277 997
rect -36 -11 89 96
<< gv2 >>
rect 47 971 49 973
rect 59 971 61 973
rect 71 971 73 973
rect 83 971 85 973
rect 95 971 97 973
rect 107 971 109 973
rect 119 971 121 973
rect 131 971 133 973
rect 143 971 145 973
rect 155 971 157 973
rect 167 971 169 973
rect 179 971 181 973
rect 191 971 193 973
rect 203 971 205 973
rect 215 971 217 973
rect 227 971 229 973
rect 239 971 241 973
rect 251 971 253 973
rect 47 959 49 961
rect 59 959 61 961
rect 71 959 73 961
rect 83 959 85 961
rect 95 959 97 961
rect 107 959 109 961
rect 119 959 121 961
rect 131 959 133 961
rect 143 959 145 961
rect 155 959 157 961
rect 167 959 169 961
rect 179 959 181 961
rect 191 959 193 961
rect 203 959 205 961
rect 215 959 217 961
rect 227 959 229 961
rect 239 959 241 961
rect 251 959 253 961
rect 47 947 49 949
rect 59 947 61 949
rect 71 947 73 949
rect 83 947 85 949
rect 95 947 97 949
rect 107 947 109 949
rect 119 947 121 949
rect 131 947 133 949
rect 143 947 145 949
rect 155 947 157 949
rect 167 947 169 949
rect 179 947 181 949
rect 191 947 193 949
rect 203 947 205 949
rect 215 947 217 949
rect 227 947 229 949
rect 239 947 241 949
rect 251 947 253 949
rect 47 935 49 937
rect 59 935 61 937
rect 71 935 73 937
rect 83 935 85 937
rect 95 935 97 937
rect 107 935 109 937
rect 119 935 121 937
rect 131 935 133 937
rect 143 935 145 937
rect 155 935 157 937
rect 167 935 169 937
rect 179 935 181 937
rect 191 935 193 937
rect 203 935 205 937
rect 215 935 217 937
rect 227 935 229 937
rect 239 935 241 937
rect 251 935 253 937
rect 47 923 49 925
rect 59 923 61 925
rect 71 923 73 925
rect 83 923 85 925
rect 95 923 97 925
rect 107 923 109 925
rect 119 923 121 925
rect 131 923 133 925
rect 143 923 145 925
rect 155 923 157 925
rect 167 923 169 925
rect 179 923 181 925
rect 191 923 193 925
rect 203 923 205 925
rect 215 923 217 925
rect 227 923 229 925
rect 239 923 241 925
rect 251 923 253 925
rect 47 911 49 913
rect 59 911 61 913
rect 71 911 73 913
rect 83 911 85 913
rect 95 911 97 913
rect 107 911 109 913
rect 119 911 121 913
rect 131 911 133 913
rect 143 911 145 913
rect 155 911 157 913
rect 167 911 169 913
rect 179 911 181 913
rect 191 911 193 913
rect 203 911 205 913
rect 215 911 217 913
rect 227 911 229 913
rect 239 911 241 913
rect 251 911 253 913
rect 47 899 49 901
rect 59 899 61 901
rect 71 899 73 901
rect 83 899 85 901
rect 95 899 97 901
rect 107 899 109 901
rect 119 899 121 901
rect 131 899 133 901
rect 143 899 145 901
rect 155 899 157 901
rect 167 899 169 901
rect 179 899 181 901
rect 191 899 193 901
rect 203 899 205 901
rect 215 899 217 901
rect 227 899 229 901
rect 239 899 241 901
rect 251 899 253 901
rect 47 887 49 889
rect 59 887 61 889
rect 71 887 73 889
rect 83 887 85 889
rect 95 887 97 889
rect 107 887 109 889
rect 119 887 121 889
rect 131 887 133 889
rect 143 887 145 889
rect 155 887 157 889
rect 167 887 169 889
rect 179 887 181 889
rect 191 887 193 889
rect 203 887 205 889
rect 215 887 217 889
rect 227 887 229 889
rect 239 887 241 889
rect 251 887 253 889
rect 47 875 49 877
rect 59 875 61 877
rect 71 875 73 877
rect 83 875 85 877
rect 95 875 97 877
rect 107 875 109 877
rect 119 875 121 877
rect 131 875 133 877
rect 143 875 145 877
rect 155 875 157 877
rect 167 875 169 877
rect 179 875 181 877
rect 191 875 193 877
rect 203 875 205 877
rect 215 875 217 877
rect 227 875 229 877
rect 239 875 241 877
rect 251 875 253 877
rect 47 863 49 865
rect 59 863 61 865
rect 71 863 73 865
rect 83 863 85 865
rect 95 863 97 865
rect 107 863 109 865
rect 119 863 121 865
rect 131 863 133 865
rect 143 863 145 865
rect 155 863 157 865
rect 167 863 169 865
rect 179 863 181 865
rect 191 863 193 865
rect 203 863 205 865
rect 215 863 217 865
rect 227 863 229 865
rect 239 863 241 865
rect 251 863 253 865
rect 47 851 49 853
rect 59 851 61 853
rect 71 851 73 853
rect 83 851 85 853
rect 95 851 97 853
rect 107 851 109 853
rect 119 851 121 853
rect 131 851 133 853
rect 143 851 145 853
rect 155 851 157 853
rect 167 851 169 853
rect 179 851 181 853
rect 191 851 193 853
rect 203 851 205 853
rect 215 851 217 853
rect 227 851 229 853
rect 239 851 241 853
rect 251 851 253 853
rect 47 839 49 841
rect 59 839 61 841
rect 71 839 73 841
rect 83 839 85 841
rect 95 839 97 841
rect 107 839 109 841
rect 119 839 121 841
rect 131 839 133 841
rect 143 839 145 841
rect 155 839 157 841
rect 167 839 169 841
rect 179 839 181 841
rect 191 839 193 841
rect 203 839 205 841
rect 215 839 217 841
rect 227 839 229 841
rect 239 839 241 841
rect 251 839 253 841
rect 47 827 49 829
rect 59 827 61 829
rect 71 827 73 829
rect 83 827 85 829
rect 95 827 97 829
rect 107 827 109 829
rect 119 827 121 829
rect 131 827 133 829
rect 143 827 145 829
rect 155 827 157 829
rect 167 827 169 829
rect 179 827 181 829
rect 191 827 193 829
rect 203 827 205 829
rect 215 827 217 829
rect 227 827 229 829
rect 239 827 241 829
rect 251 827 253 829
rect 47 815 49 817
rect 59 815 61 817
rect 71 815 73 817
rect 83 815 85 817
rect 95 815 97 817
rect 107 815 109 817
rect 119 815 121 817
rect 131 815 133 817
rect 143 815 145 817
rect 155 815 157 817
rect 167 815 169 817
rect 179 815 181 817
rect 191 815 193 817
rect 203 815 205 817
rect 215 815 217 817
rect 227 815 229 817
rect 239 815 241 817
rect 251 815 253 817
rect 47 803 49 805
rect 59 803 61 805
rect 71 803 73 805
rect 83 803 85 805
rect 95 803 97 805
rect 107 803 109 805
rect 119 803 121 805
rect 131 803 133 805
rect 143 803 145 805
rect 155 803 157 805
rect 167 803 169 805
rect 179 803 181 805
rect 191 803 193 805
rect 203 803 205 805
rect 215 803 217 805
rect 227 803 229 805
rect 239 803 241 805
rect 251 803 253 805
rect 47 791 49 793
rect 59 791 61 793
rect 71 791 73 793
rect 83 791 85 793
rect 95 791 97 793
rect 107 791 109 793
rect 119 791 121 793
rect 131 791 133 793
rect 143 791 145 793
rect 155 791 157 793
rect 167 791 169 793
rect 179 791 181 793
rect 191 791 193 793
rect 203 791 205 793
rect 215 791 217 793
rect 227 791 229 793
rect 239 791 241 793
rect 251 791 253 793
rect 47 779 49 781
rect 59 779 61 781
rect 71 779 73 781
rect 83 779 85 781
rect 95 779 97 781
rect 107 779 109 781
rect 119 779 121 781
rect 131 779 133 781
rect 143 779 145 781
rect 155 779 157 781
rect 167 779 169 781
rect 179 779 181 781
rect 191 779 193 781
rect 203 779 205 781
rect 215 779 217 781
rect 227 779 229 781
rect 239 779 241 781
rect 251 779 253 781
rect 47 767 49 769
rect 59 767 61 769
rect 71 767 73 769
rect 83 767 85 769
rect 95 767 97 769
rect 107 767 109 769
rect 119 767 121 769
rect 131 767 133 769
rect 143 767 145 769
rect 155 767 157 769
rect 167 767 169 769
rect 179 767 181 769
rect 191 767 193 769
rect 203 767 205 769
rect 215 767 217 769
rect 227 767 229 769
rect 239 767 241 769
rect 251 767 253 769
<< glass >>
rect 43 763 257 977
<< pseudo_rpoly >>
rect 126 405 191 407
rect 210 405 274 407
rect 126 393 191 395
rect 210 393 274 395
<< rpoly >>
rect 126 395 191 405
rect 210 395 274 405
<< xp >>
rect 23 743 277 997
<< labels >>
rlabel metal2 48 0 48 0 8 DO
rlabel metal2 150 0 150 0 8 DATA
rlabel metal2 261 0 261 0 8 DI
rlabel metal2 248 0 248 0 8 DIB
rlabel metal2 48 0 48 0 8 DO
rlabel metal2 15 0 15 0 8 OEN
rlabel metal2 169 129 169 129 6 gnd:2
rlabel metal2 132 535 132 535 6 vdd:2
rlabel metal2 174 307 174 307 6 Vdd!
rlabel metal2 171 364 171 364 6 Gnd!
rlabel metal1 201 404 201 404 6 hack
rlabel metal1 201 399 201 399 6 hack
rlabel metal2 48 -18 48 -18 8 DO
rlabel metal2 261 -18 261 -18 8 DI
rlabel metal2 248 -18 248 -18 8 DIB
rlabel metal2 26 -18 26 -18 8 OEN
rlabel metal1 113 -9 113 -9 8 Vdd!
rlabel metal2 97 -9 97 -9 8 GND!
<< end >>
