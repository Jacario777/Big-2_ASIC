magic
tech scmos
timestamp 1681620392
<< nwell >>
rect -8 48 32 105
<< ntransistor >>
rect 7 6 9 26
rect 12 6 14 26
<< ptransistor >>
rect 7 74 9 94
rect 15 74 17 94
<< ndiffusion >>
rect 2 6 7 26
rect 9 6 12 26
rect 14 6 19 26
<< pdiffusion >>
rect 2 74 7 94
rect 9 74 15 94
rect 17 74 22 94
<< psubstratepdiff >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratendiff >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 7 33 9 74
rect 2 29 9 33
rect 15 61 17 74
rect 15 57 22 61
rect 15 29 17 57
rect 7 26 9 29
rect 12 27 17 29
rect 12 26 14 27
rect 7 4 9 6
rect 12 4 14 6
<< genericcontact >>
rect -1 99 1 101
rect 15 99 17 101
rect 3 90 5 92
rect 11 90 13 92
rect 19 90 21 92
rect 3 85 5 87
rect 11 85 13 87
rect 19 85 21 87
rect 3 80 5 82
rect 11 80 13 82
rect 19 80 21 82
rect 3 75 5 77
rect 11 75 13 77
rect 19 75 21 77
rect 19 58 21 60
rect 3 30 5 32
rect 3 22 5 24
rect 16 22 18 24
rect 3 17 5 19
rect 16 17 18 19
rect 3 12 5 14
rect 16 12 18 14
rect 3 7 5 9
rect 16 7 18 9
rect -1 -1 1 1
rect 15 -1 17 1
<< metal1 >>
rect -2 97 26 103
rect 2 74 6 97
rect 2 29 6 37
rect 10 26 14 94
rect 18 74 22 97
rect 18 53 22 61
rect 2 3 6 26
rect 10 23 19 26
rect 15 6 19 23
rect -2 -3 26 3
<< m1p >>
rect 18 53 22 57
rect 10 43 14 47
rect 2 33 6 37
<< labels >>
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 12 45 12 45 6 Y
rlabel metal1 4 0 4 0 8 gnd
rlabel metal1 4 35 4 35 6 A
rlabel metal1 20 55 20 55 6 B
<< end >>
