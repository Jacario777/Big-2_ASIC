magic
tech scmos
timestamp 1681620392
<< nwell >>
rect 20 740 280 1000
rect 17 429 283 653
rect -3 248 303 330
rect -3 10 11 248
rect 289 10 303 248
rect -3 -4 303 10
<< ntransistor >>
rect 38 215 138 218
rect 38 170 138 173
rect 38 149 138 152
rect 38 105 138 108
rect 38 84 138 87
rect 38 40 138 43
rect 162 215 262 218
rect 162 170 262 173
rect 162 149 262 152
rect 162 105 262 108
rect 162 84 262 87
rect 162 40 262 43
<< ndiffusion >>
rect 38 218 138 227
rect 38 173 138 215
rect 38 152 138 170
rect 38 108 138 149
rect 38 87 138 105
rect 38 43 138 84
rect 38 31 138 40
rect 162 218 262 227
rect 162 173 262 215
rect 162 152 262 170
rect 162 108 262 149
rect 162 87 262 105
rect 162 43 262 84
rect 162 31 262 40
<< psubstratepdiff >>
rect 0 659 300 670
rect 0 423 11 659
rect 289 423 300 659
rect 0 343 300 423
rect 14 229 286 245
rect 14 29 30 229
rect 38 227 138 229
rect 38 29 138 31
rect 142 29 158 229
rect 162 227 262 229
rect 162 29 262 31
rect 270 29 286 229
rect 14 13 286 29
<< nsubstratendiff >>
rect 20 432 280 650
rect 0 251 300 327
rect 0 7 8 251
rect 292 7 300 251
rect 0 -1 300 7
<< polysilicon >>
rect 6 713 21 716
rect 24 713 39 716
rect 12 701 15 713
rect 24 710 27 713
rect 36 710 39 713
rect 24 707 39 710
rect 24 701 27 707
rect 36 701 39 707
rect 42 713 45 716
rect 42 710 51 713
rect 42 701 45 710
rect 48 707 51 710
rect 54 707 57 716
rect 48 704 57 707
rect 54 701 57 704
rect 60 713 63 716
rect 60 710 69 713
rect 60 701 63 710
rect 66 707 69 710
rect 72 707 75 716
rect 66 704 75 707
rect 72 701 75 704
rect 78 713 93 716
rect 96 713 111 716
rect 78 710 81 713
rect 96 710 99 713
rect 108 710 111 713
rect 78 707 93 710
rect 96 707 111 710
rect 190 707 205 710
rect 78 704 81 707
rect 78 701 93 704
rect 96 701 99 707
rect 105 701 108 707
rect 190 695 193 707
rect 196 701 199 707
rect 202 695 205 707
rect 208 707 223 710
rect 208 698 211 707
rect 220 698 223 707
rect 226 707 241 710
rect 244 707 259 710
rect 262 707 277 710
rect 226 704 229 707
rect 226 701 241 704
rect 238 698 241 701
rect 250 698 253 707
rect 262 704 265 707
rect 262 701 277 704
rect 274 698 277 701
rect 208 695 223 698
rect 226 695 241 698
rect 244 695 259 698
rect 262 695 277 698
rect 51 688 66 691
rect 69 688 84 691
rect 87 688 102 691
rect 51 679 54 688
rect 69 685 72 688
rect 87 685 90 688
rect 69 682 84 685
rect 87 682 102 685
rect 69 679 72 682
rect 99 679 102 682
rect 51 676 66 679
rect 69 676 84 679
rect 87 676 102 679
rect 31 215 38 218
rect 138 215 140 218
rect 31 173 37 215
rect 31 170 38 173
rect 138 170 140 173
rect 31 152 37 170
rect 31 149 38 152
rect 138 149 140 152
rect 31 108 37 149
rect 31 105 38 108
rect 138 105 140 108
rect 31 87 37 105
rect 31 84 38 87
rect 138 84 140 87
rect 31 43 37 84
rect 31 40 38 43
rect 138 40 140 43
rect 160 215 162 218
rect 262 215 269 218
rect 263 173 269 215
rect 160 170 162 173
rect 262 170 269 173
rect 263 152 269 170
rect 160 149 162 152
rect 262 149 269 152
rect 263 108 269 149
rect 160 105 162 108
rect 262 105 269 108
rect 263 87 269 105
rect 160 84 162 87
rect 262 84 269 87
rect 263 43 269 84
rect 160 40 162 43
rect 262 40 269 43
<< genericcontact >>
rect 2 666 4 668
rect 7 666 9 668
rect 12 666 14 668
rect 17 666 19 668
rect 22 666 24 668
rect 27 666 29 668
rect 32 666 34 668
rect 37 666 39 668
rect 42 666 44 668
rect 47 666 49 668
rect 52 666 54 668
rect 57 666 59 668
rect 62 666 64 668
rect 67 666 69 668
rect 72 666 74 668
rect 77 666 79 668
rect 82 666 84 668
rect 87 666 89 668
rect 92 666 94 668
rect 205 666 207 668
rect 210 666 212 668
rect 215 666 217 668
rect 220 666 222 668
rect 225 666 227 668
rect 230 666 232 668
rect 235 666 237 668
rect 240 666 242 668
rect 245 666 247 668
rect 250 666 252 668
rect 255 666 257 668
rect 260 666 262 668
rect 265 666 267 668
rect 270 666 272 668
rect 275 666 277 668
rect 280 666 282 668
rect 285 666 287 668
rect 290 666 292 668
rect 295 666 297 668
rect 2 661 4 663
rect 7 661 9 663
rect 12 661 14 663
rect 17 661 19 663
rect 22 661 24 663
rect 27 661 29 663
rect 32 661 34 663
rect 37 661 39 663
rect 42 661 44 663
rect 47 661 49 663
rect 52 661 54 663
rect 57 661 59 663
rect 62 661 64 663
rect 67 661 69 663
rect 72 661 74 663
rect 77 661 79 663
rect 82 661 84 663
rect 87 661 89 663
rect 92 661 94 663
rect 205 661 207 663
rect 210 661 212 663
rect 215 661 217 663
rect 220 661 222 663
rect 225 661 227 663
rect 230 661 232 663
rect 235 661 237 663
rect 240 661 242 663
rect 245 661 247 663
rect 250 661 252 663
rect 255 661 257 663
rect 260 661 262 663
rect 265 661 267 663
rect 270 661 272 663
rect 275 661 277 663
rect 280 661 282 663
rect 285 661 287 663
rect 290 661 292 663
rect 295 661 297 663
rect 2 655 4 657
rect 7 655 9 657
rect 291 655 293 657
rect 296 655 298 657
rect 2 650 4 652
rect 7 650 9 652
rect 291 650 293 652
rect 296 650 298 652
rect 2 645 4 647
rect 7 645 9 647
rect 24 646 26 648
rect 29 646 31 648
rect 34 646 36 648
rect 39 646 41 648
rect 44 646 46 648
rect 49 646 51 648
rect 54 646 56 648
rect 59 646 61 648
rect 64 646 66 648
rect 69 646 71 648
rect 74 646 76 648
rect 79 646 81 648
rect 84 646 86 648
rect 89 646 91 648
rect 94 646 96 648
rect 99 646 101 648
rect 104 646 106 648
rect 109 646 111 648
rect 114 646 116 648
rect 119 646 121 648
rect 124 646 126 648
rect 129 646 131 648
rect 134 646 136 648
rect 139 646 141 648
rect 144 646 146 648
rect 149 646 151 648
rect 154 646 156 648
rect 159 646 161 648
rect 164 646 166 648
rect 169 646 171 648
rect 174 646 176 648
rect 179 646 181 648
rect 184 646 186 648
rect 189 646 191 648
rect 194 646 196 648
rect 199 646 201 648
rect 204 646 206 648
rect 209 646 211 648
rect 214 646 216 648
rect 219 646 221 648
rect 224 646 226 648
rect 229 646 231 648
rect 234 646 236 648
rect 239 646 241 648
rect 244 646 246 648
rect 249 646 251 648
rect 254 646 256 648
rect 259 646 261 648
rect 264 646 266 648
rect 269 646 271 648
rect 274 646 276 648
rect 291 645 293 647
rect 296 645 298 647
rect 2 640 4 642
rect 7 640 9 642
rect 291 640 293 642
rect 296 640 298 642
rect 2 635 4 637
rect 7 635 9 637
rect 24 636 26 638
rect 29 636 31 638
rect 34 636 36 638
rect 39 636 41 638
rect 44 636 46 638
rect 49 636 51 638
rect 54 636 56 638
rect 59 636 61 638
rect 64 636 66 638
rect 69 636 71 638
rect 74 636 76 638
rect 79 636 81 638
rect 84 636 86 638
rect 89 636 91 638
rect 94 636 96 638
rect 99 636 101 638
rect 104 636 106 638
rect 109 636 111 638
rect 114 636 116 638
rect 119 636 121 638
rect 124 636 126 638
rect 129 636 131 638
rect 134 636 136 638
rect 139 636 141 638
rect 144 636 146 638
rect 149 636 151 638
rect 154 636 156 638
rect 159 636 161 638
rect 164 636 166 638
rect 169 636 171 638
rect 174 636 176 638
rect 179 636 181 638
rect 184 636 186 638
rect 189 636 191 638
rect 194 636 196 638
rect 199 636 201 638
rect 204 636 206 638
rect 209 636 211 638
rect 214 636 216 638
rect 219 636 221 638
rect 224 636 226 638
rect 229 636 231 638
rect 234 636 236 638
rect 239 636 241 638
rect 244 636 246 638
rect 249 636 251 638
rect 254 636 256 638
rect 259 636 261 638
rect 264 636 266 638
rect 269 636 271 638
rect 274 636 276 638
rect 291 635 293 637
rect 296 635 298 637
rect 2 630 4 632
rect 7 630 9 632
rect 291 630 293 632
rect 296 630 298 632
rect 2 625 4 627
rect 7 625 9 627
rect 24 626 26 628
rect 29 626 31 628
rect 34 626 36 628
rect 39 626 41 628
rect 44 626 46 628
rect 49 626 51 628
rect 54 626 56 628
rect 59 626 61 628
rect 64 626 66 628
rect 69 626 71 628
rect 74 626 76 628
rect 79 626 81 628
rect 84 626 86 628
rect 89 626 91 628
rect 94 626 96 628
rect 99 626 101 628
rect 104 626 106 628
rect 109 626 111 628
rect 114 626 116 628
rect 119 626 121 628
rect 124 626 126 628
rect 129 626 131 628
rect 134 626 136 628
rect 139 626 141 628
rect 144 626 146 628
rect 149 626 151 628
rect 154 626 156 628
rect 159 626 161 628
rect 164 626 166 628
rect 169 626 171 628
rect 174 626 176 628
rect 179 626 181 628
rect 184 626 186 628
rect 189 626 191 628
rect 194 626 196 628
rect 199 626 201 628
rect 204 626 206 628
rect 209 626 211 628
rect 214 626 216 628
rect 219 626 221 628
rect 224 626 226 628
rect 229 626 231 628
rect 234 626 236 628
rect 239 626 241 628
rect 244 626 246 628
rect 249 626 251 628
rect 254 626 256 628
rect 259 626 261 628
rect 264 626 266 628
rect 269 626 271 628
rect 274 626 276 628
rect 291 625 293 627
rect 296 625 298 627
rect 2 620 4 622
rect 7 620 9 622
rect 291 620 293 622
rect 296 620 298 622
rect 2 615 4 617
rect 7 615 9 617
rect 24 616 26 618
rect 29 616 31 618
rect 34 616 36 618
rect 39 616 41 618
rect 44 616 46 618
rect 49 616 51 618
rect 54 616 56 618
rect 59 616 61 618
rect 64 616 66 618
rect 69 616 71 618
rect 74 616 76 618
rect 79 616 81 618
rect 84 616 86 618
rect 89 616 91 618
rect 94 616 96 618
rect 99 616 101 618
rect 104 616 106 618
rect 109 616 111 618
rect 114 616 116 618
rect 119 616 121 618
rect 124 616 126 618
rect 129 616 131 618
rect 134 616 136 618
rect 139 616 141 618
rect 144 616 146 618
rect 149 616 151 618
rect 154 616 156 618
rect 159 616 161 618
rect 164 616 166 618
rect 169 616 171 618
rect 174 616 176 618
rect 179 616 181 618
rect 184 616 186 618
rect 189 616 191 618
rect 194 616 196 618
rect 199 616 201 618
rect 204 616 206 618
rect 209 616 211 618
rect 214 616 216 618
rect 219 616 221 618
rect 224 616 226 618
rect 229 616 231 618
rect 234 616 236 618
rect 239 616 241 618
rect 244 616 246 618
rect 249 616 251 618
rect 254 616 256 618
rect 259 616 261 618
rect 264 616 266 618
rect 269 616 271 618
rect 274 616 276 618
rect 291 615 293 617
rect 296 615 298 617
rect 2 610 4 612
rect 7 610 9 612
rect 291 610 293 612
rect 296 610 298 612
rect 2 605 4 607
rect 7 605 9 607
rect 24 606 26 608
rect 29 606 31 608
rect 34 606 36 608
rect 39 606 41 608
rect 44 606 46 608
rect 49 606 51 608
rect 54 606 56 608
rect 59 606 61 608
rect 64 606 66 608
rect 69 606 71 608
rect 74 606 76 608
rect 79 606 81 608
rect 84 606 86 608
rect 89 606 91 608
rect 94 606 96 608
rect 99 606 101 608
rect 104 606 106 608
rect 109 606 111 608
rect 114 606 116 608
rect 119 606 121 608
rect 124 606 126 608
rect 129 606 131 608
rect 134 606 136 608
rect 139 606 141 608
rect 144 606 146 608
rect 149 606 151 608
rect 154 606 156 608
rect 159 606 161 608
rect 164 606 166 608
rect 169 606 171 608
rect 174 606 176 608
rect 179 606 181 608
rect 184 606 186 608
rect 189 606 191 608
rect 194 606 196 608
rect 199 606 201 608
rect 204 606 206 608
rect 209 606 211 608
rect 214 606 216 608
rect 219 606 221 608
rect 224 606 226 608
rect 229 606 231 608
rect 234 606 236 608
rect 239 606 241 608
rect 244 606 246 608
rect 249 606 251 608
rect 254 606 256 608
rect 259 606 261 608
rect 264 606 266 608
rect 269 606 271 608
rect 274 606 276 608
rect 291 605 293 607
rect 296 605 298 607
rect 2 600 4 602
rect 7 600 9 602
rect 291 600 293 602
rect 296 600 298 602
rect 2 595 4 597
rect 7 595 9 597
rect 24 596 26 598
rect 29 596 31 598
rect 34 596 36 598
rect 39 596 41 598
rect 44 596 46 598
rect 49 596 51 598
rect 54 596 56 598
rect 59 596 61 598
rect 64 596 66 598
rect 69 596 71 598
rect 74 596 76 598
rect 79 596 81 598
rect 84 596 86 598
rect 89 596 91 598
rect 94 596 96 598
rect 99 596 101 598
rect 104 596 106 598
rect 109 596 111 598
rect 114 596 116 598
rect 119 596 121 598
rect 124 596 126 598
rect 129 596 131 598
rect 134 596 136 598
rect 139 596 141 598
rect 144 596 146 598
rect 149 596 151 598
rect 154 596 156 598
rect 159 596 161 598
rect 164 596 166 598
rect 169 596 171 598
rect 174 596 176 598
rect 179 596 181 598
rect 184 596 186 598
rect 189 596 191 598
rect 194 596 196 598
rect 199 596 201 598
rect 204 596 206 598
rect 209 596 211 598
rect 214 596 216 598
rect 219 596 221 598
rect 224 596 226 598
rect 229 596 231 598
rect 234 596 236 598
rect 239 596 241 598
rect 244 596 246 598
rect 249 596 251 598
rect 254 596 256 598
rect 259 596 261 598
rect 264 596 266 598
rect 269 596 271 598
rect 274 596 276 598
rect 291 595 293 597
rect 296 595 298 597
rect 2 590 4 592
rect 7 590 9 592
rect 291 590 293 592
rect 296 590 298 592
rect 2 585 4 587
rect 7 585 9 587
rect 24 586 26 588
rect 29 586 31 588
rect 34 586 36 588
rect 39 586 41 588
rect 44 586 46 588
rect 49 586 51 588
rect 54 586 56 588
rect 59 586 61 588
rect 64 586 66 588
rect 69 586 71 588
rect 74 586 76 588
rect 79 586 81 588
rect 84 586 86 588
rect 89 586 91 588
rect 94 586 96 588
rect 99 586 101 588
rect 104 586 106 588
rect 109 586 111 588
rect 114 586 116 588
rect 119 586 121 588
rect 124 586 126 588
rect 129 586 131 588
rect 134 586 136 588
rect 139 586 141 588
rect 144 586 146 588
rect 149 586 151 588
rect 154 586 156 588
rect 159 586 161 588
rect 164 586 166 588
rect 169 586 171 588
rect 174 586 176 588
rect 179 586 181 588
rect 184 586 186 588
rect 189 586 191 588
rect 194 586 196 588
rect 199 586 201 588
rect 204 586 206 588
rect 209 586 211 588
rect 214 586 216 588
rect 219 586 221 588
rect 224 586 226 588
rect 229 586 231 588
rect 234 586 236 588
rect 239 586 241 588
rect 244 586 246 588
rect 249 586 251 588
rect 254 586 256 588
rect 259 586 261 588
rect 264 586 266 588
rect 269 586 271 588
rect 274 586 276 588
rect 291 585 293 587
rect 296 585 298 587
rect 2 580 4 582
rect 7 580 9 582
rect 291 580 293 582
rect 296 580 298 582
rect 2 575 4 577
rect 7 575 9 577
rect 24 576 26 578
rect 29 576 31 578
rect 34 576 36 578
rect 39 576 41 578
rect 44 576 46 578
rect 49 576 51 578
rect 54 576 56 578
rect 59 576 61 578
rect 64 576 66 578
rect 69 576 71 578
rect 74 576 76 578
rect 79 576 81 578
rect 84 576 86 578
rect 89 576 91 578
rect 94 576 96 578
rect 99 576 101 578
rect 104 576 106 578
rect 109 576 111 578
rect 114 576 116 578
rect 119 576 121 578
rect 124 576 126 578
rect 129 576 131 578
rect 134 576 136 578
rect 139 576 141 578
rect 144 576 146 578
rect 149 576 151 578
rect 154 576 156 578
rect 159 576 161 578
rect 164 576 166 578
rect 169 576 171 578
rect 174 576 176 578
rect 179 576 181 578
rect 184 576 186 578
rect 189 576 191 578
rect 194 576 196 578
rect 199 576 201 578
rect 204 576 206 578
rect 209 576 211 578
rect 214 576 216 578
rect 219 576 221 578
rect 224 576 226 578
rect 229 576 231 578
rect 234 576 236 578
rect 239 576 241 578
rect 244 576 246 578
rect 249 576 251 578
rect 254 576 256 578
rect 259 576 261 578
rect 264 576 266 578
rect 269 576 271 578
rect 274 576 276 578
rect 291 575 293 577
rect 296 575 298 577
rect 2 570 4 572
rect 7 570 9 572
rect 291 570 293 572
rect 296 570 298 572
rect 2 565 4 567
rect 7 565 9 567
rect 24 566 26 568
rect 29 566 31 568
rect 34 566 36 568
rect 39 566 41 568
rect 44 566 46 568
rect 49 566 51 568
rect 54 566 56 568
rect 59 566 61 568
rect 64 566 66 568
rect 69 566 71 568
rect 74 566 76 568
rect 79 566 81 568
rect 84 566 86 568
rect 89 566 91 568
rect 94 566 96 568
rect 99 566 101 568
rect 104 566 106 568
rect 109 566 111 568
rect 114 566 116 568
rect 119 566 121 568
rect 124 566 126 568
rect 129 566 131 568
rect 134 566 136 568
rect 139 566 141 568
rect 144 566 146 568
rect 149 566 151 568
rect 154 566 156 568
rect 159 566 161 568
rect 164 566 166 568
rect 169 566 171 568
rect 174 566 176 568
rect 179 566 181 568
rect 184 566 186 568
rect 189 566 191 568
rect 194 566 196 568
rect 199 566 201 568
rect 204 566 206 568
rect 209 566 211 568
rect 214 566 216 568
rect 219 566 221 568
rect 224 566 226 568
rect 229 566 231 568
rect 234 566 236 568
rect 239 566 241 568
rect 244 566 246 568
rect 249 566 251 568
rect 254 566 256 568
rect 259 566 261 568
rect 264 566 266 568
rect 269 566 271 568
rect 274 566 276 568
rect 291 565 293 567
rect 296 565 298 567
rect 2 560 4 562
rect 7 560 9 562
rect 291 560 293 562
rect 296 560 298 562
rect 2 555 4 557
rect 7 555 9 557
rect 24 556 26 558
rect 29 556 31 558
rect 34 556 36 558
rect 39 556 41 558
rect 44 556 46 558
rect 49 556 51 558
rect 54 556 56 558
rect 59 556 61 558
rect 64 556 66 558
rect 69 556 71 558
rect 74 556 76 558
rect 79 556 81 558
rect 84 556 86 558
rect 89 556 91 558
rect 94 556 96 558
rect 99 556 101 558
rect 104 556 106 558
rect 109 556 111 558
rect 114 556 116 558
rect 119 556 121 558
rect 124 556 126 558
rect 129 556 131 558
rect 134 556 136 558
rect 139 556 141 558
rect 144 556 146 558
rect 149 556 151 558
rect 154 556 156 558
rect 159 556 161 558
rect 164 556 166 558
rect 169 556 171 558
rect 174 556 176 558
rect 179 556 181 558
rect 184 556 186 558
rect 189 556 191 558
rect 194 556 196 558
rect 199 556 201 558
rect 204 556 206 558
rect 209 556 211 558
rect 214 556 216 558
rect 219 556 221 558
rect 224 556 226 558
rect 229 556 231 558
rect 234 556 236 558
rect 239 556 241 558
rect 244 556 246 558
rect 249 556 251 558
rect 254 556 256 558
rect 259 556 261 558
rect 264 556 266 558
rect 269 556 271 558
rect 274 556 276 558
rect 291 555 293 557
rect 296 555 298 557
rect 2 550 4 552
rect 7 550 9 552
rect 291 550 293 552
rect 296 550 298 552
rect 2 545 4 547
rect 7 545 9 547
rect 24 546 26 548
rect 29 546 31 548
rect 34 546 36 548
rect 39 546 41 548
rect 44 546 46 548
rect 49 546 51 548
rect 54 546 56 548
rect 59 546 61 548
rect 64 546 66 548
rect 69 546 71 548
rect 74 546 76 548
rect 79 546 81 548
rect 84 546 86 548
rect 89 546 91 548
rect 94 546 96 548
rect 99 546 101 548
rect 104 546 106 548
rect 109 546 111 548
rect 114 546 116 548
rect 119 546 121 548
rect 124 546 126 548
rect 129 546 131 548
rect 134 546 136 548
rect 139 546 141 548
rect 144 546 146 548
rect 149 546 151 548
rect 154 546 156 548
rect 159 546 161 548
rect 164 546 166 548
rect 169 546 171 548
rect 174 546 176 548
rect 179 546 181 548
rect 184 546 186 548
rect 189 546 191 548
rect 194 546 196 548
rect 199 546 201 548
rect 204 546 206 548
rect 209 546 211 548
rect 214 546 216 548
rect 219 546 221 548
rect 224 546 226 548
rect 229 546 231 548
rect 234 546 236 548
rect 239 546 241 548
rect 244 546 246 548
rect 249 546 251 548
rect 254 546 256 548
rect 259 546 261 548
rect 264 546 266 548
rect 269 546 271 548
rect 274 546 276 548
rect 291 545 293 547
rect 296 545 298 547
rect 2 540 4 542
rect 7 540 9 542
rect 291 540 293 542
rect 296 540 298 542
rect 2 535 4 537
rect 7 535 9 537
rect 24 536 26 538
rect 29 536 31 538
rect 34 536 36 538
rect 39 536 41 538
rect 44 536 46 538
rect 49 536 51 538
rect 54 536 56 538
rect 59 536 61 538
rect 64 536 66 538
rect 69 536 71 538
rect 74 536 76 538
rect 79 536 81 538
rect 84 536 86 538
rect 89 536 91 538
rect 94 536 96 538
rect 99 536 101 538
rect 104 536 106 538
rect 109 536 111 538
rect 114 536 116 538
rect 119 536 121 538
rect 124 536 126 538
rect 129 536 131 538
rect 134 536 136 538
rect 139 536 141 538
rect 144 536 146 538
rect 149 536 151 538
rect 154 536 156 538
rect 159 536 161 538
rect 164 536 166 538
rect 169 536 171 538
rect 174 536 176 538
rect 179 536 181 538
rect 184 536 186 538
rect 189 536 191 538
rect 194 536 196 538
rect 199 536 201 538
rect 204 536 206 538
rect 209 536 211 538
rect 214 536 216 538
rect 219 536 221 538
rect 224 536 226 538
rect 229 536 231 538
rect 234 536 236 538
rect 239 536 241 538
rect 244 536 246 538
rect 249 536 251 538
rect 254 536 256 538
rect 259 536 261 538
rect 264 536 266 538
rect 269 536 271 538
rect 274 536 276 538
rect 291 535 293 537
rect 296 535 298 537
rect 2 530 4 532
rect 7 530 9 532
rect 291 530 293 532
rect 296 530 298 532
rect 2 525 4 527
rect 7 525 9 527
rect 24 526 26 528
rect 29 526 31 528
rect 34 526 36 528
rect 39 526 41 528
rect 44 526 46 528
rect 49 526 51 528
rect 54 526 56 528
rect 59 526 61 528
rect 64 526 66 528
rect 69 526 71 528
rect 74 526 76 528
rect 79 526 81 528
rect 84 526 86 528
rect 89 526 91 528
rect 94 526 96 528
rect 99 526 101 528
rect 104 526 106 528
rect 109 526 111 528
rect 114 526 116 528
rect 119 526 121 528
rect 124 526 126 528
rect 129 526 131 528
rect 134 526 136 528
rect 139 526 141 528
rect 144 526 146 528
rect 149 526 151 528
rect 154 526 156 528
rect 159 526 161 528
rect 164 526 166 528
rect 169 526 171 528
rect 174 526 176 528
rect 179 526 181 528
rect 184 526 186 528
rect 189 526 191 528
rect 194 526 196 528
rect 199 526 201 528
rect 204 526 206 528
rect 209 526 211 528
rect 214 526 216 528
rect 219 526 221 528
rect 224 526 226 528
rect 229 526 231 528
rect 234 526 236 528
rect 239 526 241 528
rect 244 526 246 528
rect 249 526 251 528
rect 254 526 256 528
rect 259 526 261 528
rect 264 526 266 528
rect 269 526 271 528
rect 274 526 276 528
rect 291 525 293 527
rect 296 525 298 527
rect 2 520 4 522
rect 7 520 9 522
rect 291 520 293 522
rect 296 520 298 522
rect 2 515 4 517
rect 7 515 9 517
rect 24 516 26 518
rect 29 516 31 518
rect 34 516 36 518
rect 39 516 41 518
rect 44 516 46 518
rect 49 516 51 518
rect 54 516 56 518
rect 59 516 61 518
rect 64 516 66 518
rect 69 516 71 518
rect 74 516 76 518
rect 79 516 81 518
rect 84 516 86 518
rect 89 516 91 518
rect 94 516 96 518
rect 99 516 101 518
rect 104 516 106 518
rect 109 516 111 518
rect 114 516 116 518
rect 119 516 121 518
rect 124 516 126 518
rect 129 516 131 518
rect 134 516 136 518
rect 139 516 141 518
rect 144 516 146 518
rect 149 516 151 518
rect 154 516 156 518
rect 159 516 161 518
rect 164 516 166 518
rect 169 516 171 518
rect 174 516 176 518
rect 179 516 181 518
rect 184 516 186 518
rect 189 516 191 518
rect 194 516 196 518
rect 199 516 201 518
rect 204 516 206 518
rect 209 516 211 518
rect 214 516 216 518
rect 219 516 221 518
rect 224 516 226 518
rect 229 516 231 518
rect 234 516 236 518
rect 239 516 241 518
rect 244 516 246 518
rect 249 516 251 518
rect 254 516 256 518
rect 259 516 261 518
rect 264 516 266 518
rect 269 516 271 518
rect 274 516 276 518
rect 291 515 293 517
rect 296 515 298 517
rect 2 510 4 512
rect 7 510 9 512
rect 291 510 293 512
rect 296 510 298 512
rect 2 505 4 507
rect 7 505 9 507
rect 24 506 26 508
rect 29 506 31 508
rect 34 506 36 508
rect 39 506 41 508
rect 44 506 46 508
rect 49 506 51 508
rect 54 506 56 508
rect 59 506 61 508
rect 64 506 66 508
rect 69 506 71 508
rect 74 506 76 508
rect 79 506 81 508
rect 84 506 86 508
rect 89 506 91 508
rect 94 506 96 508
rect 99 506 101 508
rect 104 506 106 508
rect 109 506 111 508
rect 114 506 116 508
rect 119 506 121 508
rect 124 506 126 508
rect 129 506 131 508
rect 134 506 136 508
rect 139 506 141 508
rect 144 506 146 508
rect 149 506 151 508
rect 154 506 156 508
rect 159 506 161 508
rect 164 506 166 508
rect 169 506 171 508
rect 174 506 176 508
rect 179 506 181 508
rect 184 506 186 508
rect 189 506 191 508
rect 194 506 196 508
rect 199 506 201 508
rect 204 506 206 508
rect 209 506 211 508
rect 214 506 216 508
rect 219 506 221 508
rect 224 506 226 508
rect 229 506 231 508
rect 234 506 236 508
rect 239 506 241 508
rect 244 506 246 508
rect 249 506 251 508
rect 254 506 256 508
rect 259 506 261 508
rect 264 506 266 508
rect 269 506 271 508
rect 274 506 276 508
rect 291 505 293 507
rect 296 505 298 507
rect 2 500 4 502
rect 7 500 9 502
rect 291 500 293 502
rect 296 500 298 502
rect 2 495 4 497
rect 7 495 9 497
rect 24 496 26 498
rect 29 496 31 498
rect 34 496 36 498
rect 39 496 41 498
rect 44 496 46 498
rect 49 496 51 498
rect 54 496 56 498
rect 59 496 61 498
rect 64 496 66 498
rect 69 496 71 498
rect 74 496 76 498
rect 79 496 81 498
rect 84 496 86 498
rect 89 496 91 498
rect 94 496 96 498
rect 99 496 101 498
rect 104 496 106 498
rect 109 496 111 498
rect 114 496 116 498
rect 119 496 121 498
rect 124 496 126 498
rect 129 496 131 498
rect 134 496 136 498
rect 139 496 141 498
rect 144 496 146 498
rect 149 496 151 498
rect 154 496 156 498
rect 159 496 161 498
rect 164 496 166 498
rect 169 496 171 498
rect 174 496 176 498
rect 179 496 181 498
rect 184 496 186 498
rect 189 496 191 498
rect 194 496 196 498
rect 199 496 201 498
rect 204 496 206 498
rect 209 496 211 498
rect 214 496 216 498
rect 219 496 221 498
rect 224 496 226 498
rect 229 496 231 498
rect 234 496 236 498
rect 239 496 241 498
rect 244 496 246 498
rect 249 496 251 498
rect 254 496 256 498
rect 259 496 261 498
rect 264 496 266 498
rect 269 496 271 498
rect 274 496 276 498
rect 291 495 293 497
rect 296 495 298 497
rect 2 490 4 492
rect 7 490 9 492
rect 291 490 293 492
rect 296 490 298 492
rect 2 485 4 487
rect 7 485 9 487
rect 24 486 26 488
rect 29 486 31 488
rect 34 486 36 488
rect 39 486 41 488
rect 44 486 46 488
rect 49 486 51 488
rect 54 486 56 488
rect 59 486 61 488
rect 64 486 66 488
rect 69 486 71 488
rect 74 486 76 488
rect 79 486 81 488
rect 84 486 86 488
rect 89 486 91 488
rect 94 486 96 488
rect 99 486 101 488
rect 104 486 106 488
rect 109 486 111 488
rect 114 486 116 488
rect 119 486 121 488
rect 124 486 126 488
rect 129 486 131 488
rect 134 486 136 488
rect 139 486 141 488
rect 144 486 146 488
rect 149 486 151 488
rect 154 486 156 488
rect 159 486 161 488
rect 164 486 166 488
rect 169 486 171 488
rect 174 486 176 488
rect 179 486 181 488
rect 184 486 186 488
rect 189 486 191 488
rect 194 486 196 488
rect 199 486 201 488
rect 204 486 206 488
rect 209 486 211 488
rect 214 486 216 488
rect 219 486 221 488
rect 224 486 226 488
rect 229 486 231 488
rect 234 486 236 488
rect 239 486 241 488
rect 244 486 246 488
rect 249 486 251 488
rect 254 486 256 488
rect 259 486 261 488
rect 264 486 266 488
rect 269 486 271 488
rect 274 486 276 488
rect 291 485 293 487
rect 296 485 298 487
rect 2 480 4 482
rect 7 480 9 482
rect 291 480 293 482
rect 296 480 298 482
rect 2 475 4 477
rect 7 475 9 477
rect 24 476 26 478
rect 29 476 31 478
rect 34 476 36 478
rect 39 476 41 478
rect 44 476 46 478
rect 49 476 51 478
rect 54 476 56 478
rect 59 476 61 478
rect 64 476 66 478
rect 69 476 71 478
rect 74 476 76 478
rect 79 476 81 478
rect 84 476 86 478
rect 89 476 91 478
rect 94 476 96 478
rect 99 476 101 478
rect 104 476 106 478
rect 109 476 111 478
rect 114 476 116 478
rect 119 476 121 478
rect 124 476 126 478
rect 129 476 131 478
rect 134 476 136 478
rect 139 476 141 478
rect 144 476 146 478
rect 149 476 151 478
rect 154 476 156 478
rect 159 476 161 478
rect 164 476 166 478
rect 169 476 171 478
rect 174 476 176 478
rect 179 476 181 478
rect 184 476 186 478
rect 189 476 191 478
rect 194 476 196 478
rect 199 476 201 478
rect 204 476 206 478
rect 209 476 211 478
rect 214 476 216 478
rect 219 476 221 478
rect 224 476 226 478
rect 229 476 231 478
rect 234 476 236 478
rect 239 476 241 478
rect 244 476 246 478
rect 249 476 251 478
rect 254 476 256 478
rect 259 476 261 478
rect 264 476 266 478
rect 269 476 271 478
rect 274 476 276 478
rect 291 475 293 477
rect 296 475 298 477
rect 2 470 4 472
rect 7 470 9 472
rect 291 470 293 472
rect 296 470 298 472
rect 2 465 4 467
rect 7 465 9 467
rect 24 466 26 468
rect 29 466 31 468
rect 34 466 36 468
rect 39 466 41 468
rect 44 466 46 468
rect 49 466 51 468
rect 54 466 56 468
rect 59 466 61 468
rect 64 466 66 468
rect 69 466 71 468
rect 74 466 76 468
rect 79 466 81 468
rect 84 466 86 468
rect 89 466 91 468
rect 94 466 96 468
rect 99 466 101 468
rect 104 466 106 468
rect 109 466 111 468
rect 114 466 116 468
rect 119 466 121 468
rect 124 466 126 468
rect 129 466 131 468
rect 134 466 136 468
rect 139 466 141 468
rect 144 466 146 468
rect 149 466 151 468
rect 154 466 156 468
rect 159 466 161 468
rect 164 466 166 468
rect 169 466 171 468
rect 174 466 176 468
rect 179 466 181 468
rect 184 466 186 468
rect 189 466 191 468
rect 194 466 196 468
rect 199 466 201 468
rect 204 466 206 468
rect 209 466 211 468
rect 214 466 216 468
rect 219 466 221 468
rect 224 466 226 468
rect 229 466 231 468
rect 234 466 236 468
rect 239 466 241 468
rect 244 466 246 468
rect 249 466 251 468
rect 254 466 256 468
rect 259 466 261 468
rect 264 466 266 468
rect 269 466 271 468
rect 274 466 276 468
rect 291 465 293 467
rect 296 465 298 467
rect 2 460 4 462
rect 7 460 9 462
rect 291 460 293 462
rect 296 460 298 462
rect 2 455 4 457
rect 7 455 9 457
rect 24 456 26 458
rect 29 456 31 458
rect 34 456 36 458
rect 39 456 41 458
rect 44 456 46 458
rect 49 456 51 458
rect 54 456 56 458
rect 59 456 61 458
rect 64 456 66 458
rect 69 456 71 458
rect 74 456 76 458
rect 79 456 81 458
rect 84 456 86 458
rect 89 456 91 458
rect 94 456 96 458
rect 99 456 101 458
rect 104 456 106 458
rect 109 456 111 458
rect 114 456 116 458
rect 119 456 121 458
rect 124 456 126 458
rect 129 456 131 458
rect 134 456 136 458
rect 139 456 141 458
rect 144 456 146 458
rect 149 456 151 458
rect 154 456 156 458
rect 159 456 161 458
rect 164 456 166 458
rect 169 456 171 458
rect 174 456 176 458
rect 179 456 181 458
rect 184 456 186 458
rect 189 456 191 458
rect 194 456 196 458
rect 199 456 201 458
rect 204 456 206 458
rect 209 456 211 458
rect 214 456 216 458
rect 219 456 221 458
rect 224 456 226 458
rect 229 456 231 458
rect 234 456 236 458
rect 239 456 241 458
rect 244 456 246 458
rect 249 456 251 458
rect 254 456 256 458
rect 259 456 261 458
rect 264 456 266 458
rect 269 456 271 458
rect 274 456 276 458
rect 291 455 293 457
rect 296 455 298 457
rect 2 450 4 452
rect 7 450 9 452
rect 291 450 293 452
rect 296 450 298 452
rect 2 445 4 447
rect 7 445 9 447
rect 24 446 26 448
rect 29 446 31 448
rect 34 446 36 448
rect 39 446 41 448
rect 44 446 46 448
rect 49 446 51 448
rect 54 446 56 448
rect 59 446 61 448
rect 64 446 66 448
rect 69 446 71 448
rect 74 446 76 448
rect 79 446 81 448
rect 84 446 86 448
rect 89 446 91 448
rect 94 446 96 448
rect 99 446 101 448
rect 104 446 106 448
rect 109 446 111 448
rect 114 446 116 448
rect 119 446 121 448
rect 124 446 126 448
rect 129 446 131 448
rect 134 446 136 448
rect 139 446 141 448
rect 144 446 146 448
rect 149 446 151 448
rect 154 446 156 448
rect 159 446 161 448
rect 164 446 166 448
rect 169 446 171 448
rect 174 446 176 448
rect 179 446 181 448
rect 184 446 186 448
rect 189 446 191 448
rect 194 446 196 448
rect 199 446 201 448
rect 204 446 206 448
rect 209 446 211 448
rect 214 446 216 448
rect 219 446 221 448
rect 224 446 226 448
rect 229 446 231 448
rect 234 446 236 448
rect 239 446 241 448
rect 244 446 246 448
rect 249 446 251 448
rect 254 446 256 448
rect 259 446 261 448
rect 264 446 266 448
rect 269 446 271 448
rect 274 446 276 448
rect 291 445 293 447
rect 296 445 298 447
rect 2 440 4 442
rect 7 440 9 442
rect 291 440 293 442
rect 296 440 298 442
rect 2 435 4 437
rect 7 435 9 437
rect 24 436 26 438
rect 29 436 31 438
rect 34 436 36 438
rect 39 436 41 438
rect 44 436 46 438
rect 49 436 51 438
rect 54 436 56 438
rect 59 436 61 438
rect 64 436 66 438
rect 69 436 71 438
rect 74 436 76 438
rect 79 436 81 438
rect 84 436 86 438
rect 89 436 91 438
rect 94 436 96 438
rect 99 436 101 438
rect 104 436 106 438
rect 109 436 111 438
rect 114 436 116 438
rect 119 436 121 438
rect 124 436 126 438
rect 129 436 131 438
rect 134 436 136 438
rect 139 436 141 438
rect 144 436 146 438
rect 149 436 151 438
rect 154 436 156 438
rect 159 436 161 438
rect 164 436 166 438
rect 169 436 171 438
rect 174 436 176 438
rect 179 436 181 438
rect 184 436 186 438
rect 189 436 191 438
rect 194 436 196 438
rect 199 436 201 438
rect 204 436 206 438
rect 209 436 211 438
rect 214 436 216 438
rect 219 436 221 438
rect 224 436 226 438
rect 229 436 231 438
rect 234 436 236 438
rect 239 436 241 438
rect 244 436 246 438
rect 249 436 251 438
rect 254 436 256 438
rect 259 436 261 438
rect 264 436 266 438
rect 269 436 271 438
rect 274 436 276 438
rect 291 435 293 437
rect 296 435 298 437
rect 2 430 4 432
rect 7 430 9 432
rect 291 430 293 432
rect 296 430 298 432
rect 2 425 4 427
rect 7 425 9 427
rect 291 425 293 427
rect 296 425 298 427
rect 144 415 146 417
rect 149 415 151 417
rect 154 415 156 417
rect 205 415 207 417
rect 210 415 212 417
rect 215 415 217 417
rect 220 415 222 417
rect 225 415 227 417
rect 230 415 232 417
rect 235 415 237 417
rect 240 415 242 417
rect 245 415 247 417
rect 250 415 252 417
rect 255 415 257 417
rect 260 415 262 417
rect 265 415 267 417
rect 270 415 272 417
rect 275 415 277 417
rect 280 415 282 417
rect 285 415 287 417
rect 290 415 292 417
rect 295 415 297 417
rect 3 410 5 412
rect 8 410 10 412
rect 13 410 15 412
rect 18 410 20 412
rect 23 410 25 412
rect 28 410 30 412
rect 33 410 35 412
rect 38 410 40 412
rect 43 410 45 412
rect 48 410 50 412
rect 53 410 55 412
rect 58 410 60 412
rect 63 410 65 412
rect 68 410 70 412
rect 73 410 75 412
rect 78 410 80 412
rect 83 410 85 412
rect 88 410 90 412
rect 93 410 95 412
rect 144 405 146 407
rect 149 405 151 407
rect 154 405 156 407
rect 205 405 207 407
rect 210 405 212 407
rect 215 405 217 407
rect 220 405 222 407
rect 225 405 227 407
rect 230 405 232 407
rect 235 405 237 407
rect 240 405 242 407
rect 245 405 247 407
rect 250 405 252 407
rect 255 405 257 407
rect 260 405 262 407
rect 265 405 267 407
rect 270 405 272 407
rect 275 405 277 407
rect 280 405 282 407
rect 285 405 287 407
rect 290 405 292 407
rect 295 405 297 407
rect 3 400 5 402
rect 8 400 10 402
rect 13 400 15 402
rect 18 400 20 402
rect 23 400 25 402
rect 28 400 30 402
rect 33 400 35 402
rect 38 400 40 402
rect 43 400 45 402
rect 48 400 50 402
rect 53 400 55 402
rect 58 400 60 402
rect 63 400 65 402
rect 68 400 70 402
rect 73 400 75 402
rect 78 400 80 402
rect 83 400 85 402
rect 88 400 90 402
rect 93 400 95 402
rect 144 395 146 397
rect 149 395 151 397
rect 154 395 156 397
rect 205 395 207 397
rect 210 395 212 397
rect 215 395 217 397
rect 220 395 222 397
rect 225 395 227 397
rect 230 395 232 397
rect 235 395 237 397
rect 240 395 242 397
rect 245 395 247 397
rect 250 395 252 397
rect 255 395 257 397
rect 260 395 262 397
rect 265 395 267 397
rect 270 395 272 397
rect 275 395 277 397
rect 280 395 282 397
rect 285 395 287 397
rect 290 395 292 397
rect 295 395 297 397
rect 3 390 5 392
rect 8 390 10 392
rect 13 390 15 392
rect 18 390 20 392
rect 23 390 25 392
rect 28 390 30 392
rect 33 390 35 392
rect 38 390 40 392
rect 43 390 45 392
rect 48 390 50 392
rect 53 390 55 392
rect 58 390 60 392
rect 63 390 65 392
rect 68 390 70 392
rect 73 390 75 392
rect 78 390 80 392
rect 83 390 85 392
rect 88 390 90 392
rect 93 390 95 392
rect 144 385 146 387
rect 149 385 151 387
rect 154 385 156 387
rect 205 385 207 387
rect 210 385 212 387
rect 215 385 217 387
rect 220 385 222 387
rect 225 385 227 387
rect 230 385 232 387
rect 235 385 237 387
rect 240 385 242 387
rect 245 385 247 387
rect 250 385 252 387
rect 255 385 257 387
rect 260 385 262 387
rect 265 385 267 387
rect 270 385 272 387
rect 275 385 277 387
rect 280 385 282 387
rect 285 385 287 387
rect 290 385 292 387
rect 295 385 297 387
rect 3 380 5 382
rect 8 380 10 382
rect 13 380 15 382
rect 18 380 20 382
rect 23 380 25 382
rect 28 380 30 382
rect 33 380 35 382
rect 38 380 40 382
rect 43 380 45 382
rect 48 380 50 382
rect 53 380 55 382
rect 58 380 60 382
rect 63 380 65 382
rect 68 380 70 382
rect 73 380 75 382
rect 78 380 80 382
rect 83 380 85 382
rect 88 380 90 382
rect 93 380 95 382
rect 144 375 146 377
rect 149 375 151 377
rect 154 375 156 377
rect 205 375 207 377
rect 210 375 212 377
rect 215 375 217 377
rect 220 375 222 377
rect 225 375 227 377
rect 230 375 232 377
rect 235 375 237 377
rect 240 375 242 377
rect 245 375 247 377
rect 250 375 252 377
rect 255 375 257 377
rect 260 375 262 377
rect 265 375 267 377
rect 270 375 272 377
rect 275 375 277 377
rect 280 375 282 377
rect 285 375 287 377
rect 290 375 292 377
rect 295 375 297 377
rect 3 370 5 372
rect 8 370 10 372
rect 13 370 15 372
rect 18 370 20 372
rect 23 370 25 372
rect 28 370 30 372
rect 33 370 35 372
rect 38 370 40 372
rect 43 370 45 372
rect 48 370 50 372
rect 53 370 55 372
rect 58 370 60 372
rect 63 370 65 372
rect 68 370 70 372
rect 73 370 75 372
rect 78 370 80 372
rect 83 370 85 372
rect 88 370 90 372
rect 93 370 95 372
rect 144 365 146 367
rect 149 365 151 367
rect 154 365 156 367
rect 205 365 207 367
rect 210 365 212 367
rect 215 365 217 367
rect 220 365 222 367
rect 225 365 227 367
rect 230 365 232 367
rect 235 365 237 367
rect 240 365 242 367
rect 245 365 247 367
rect 250 365 252 367
rect 255 365 257 367
rect 260 365 262 367
rect 265 365 267 367
rect 270 365 272 367
rect 275 365 277 367
rect 280 365 282 367
rect 285 365 287 367
rect 290 365 292 367
rect 295 365 297 367
rect 3 360 5 362
rect 8 360 10 362
rect 13 360 15 362
rect 18 360 20 362
rect 23 360 25 362
rect 28 360 30 362
rect 33 360 35 362
rect 38 360 40 362
rect 43 360 45 362
rect 48 360 50 362
rect 53 360 55 362
rect 58 360 60 362
rect 63 360 65 362
rect 68 360 70 362
rect 73 360 75 362
rect 78 360 80 362
rect 83 360 85 362
rect 88 360 90 362
rect 93 360 95 362
rect 144 355 146 357
rect 149 355 151 357
rect 154 355 156 357
rect 205 355 207 357
rect 210 355 212 357
rect 215 355 217 357
rect 220 355 222 357
rect 225 355 227 357
rect 230 355 232 357
rect 235 355 237 357
rect 240 355 242 357
rect 245 355 247 357
rect 250 355 252 357
rect 255 355 257 357
rect 260 355 262 357
rect 265 355 267 357
rect 270 355 272 357
rect 275 355 277 357
rect 280 355 282 357
rect 285 355 287 357
rect 290 355 292 357
rect 295 355 297 357
rect 3 345 5 347
rect 8 345 10 347
rect 13 345 15 347
rect 18 345 20 347
rect 23 345 25 347
rect 28 345 30 347
rect 33 345 35 347
rect 38 345 40 347
rect 43 345 45 347
rect 48 345 50 347
rect 53 345 55 347
rect 58 345 60 347
rect 63 345 65 347
rect 68 345 70 347
rect 73 345 75 347
rect 78 345 80 347
rect 83 345 85 347
rect 88 345 90 347
rect 93 345 95 347
rect 144 345 146 347
rect 149 345 151 347
rect 154 345 156 347
rect 205 345 207 347
rect 210 345 212 347
rect 215 345 217 347
rect 220 345 222 347
rect 225 345 227 347
rect 230 345 232 347
rect 235 345 237 347
rect 240 345 242 347
rect 245 345 247 347
rect 250 345 252 347
rect 255 345 257 347
rect 260 345 262 347
rect 265 345 267 347
rect 270 345 272 347
rect 275 345 277 347
rect 280 345 282 347
rect 285 345 287 347
rect 290 345 292 347
rect 295 345 297 347
rect 4 323 6 325
rect 9 323 11 325
rect 14 323 16 325
rect 19 323 21 325
rect 24 323 26 325
rect 29 323 31 325
rect 34 323 36 325
rect 39 323 41 325
rect 44 323 46 325
rect 49 323 51 325
rect 54 323 56 325
rect 59 323 61 325
rect 64 323 66 325
rect 69 323 71 325
rect 74 323 76 325
rect 79 323 81 325
rect 84 323 86 325
rect 89 323 91 325
rect 94 323 96 325
rect 99 323 101 325
rect 104 323 106 325
rect 109 323 111 325
rect 114 323 116 325
rect 119 323 121 325
rect 124 323 126 325
rect 129 323 131 325
rect 134 323 136 325
rect 139 323 141 325
rect 144 323 146 325
rect 149 323 151 325
rect 154 323 156 325
rect 159 323 161 325
rect 164 323 166 325
rect 169 323 171 325
rect 174 323 176 325
rect 179 323 181 325
rect 184 323 186 325
rect 189 323 191 325
rect 194 323 196 325
rect 199 323 201 325
rect 204 323 206 325
rect 209 323 211 325
rect 214 323 216 325
rect 219 323 221 325
rect 224 323 226 325
rect 229 323 231 325
rect 234 323 236 325
rect 239 323 241 325
rect 244 323 246 325
rect 249 323 251 325
rect 254 323 256 325
rect 259 323 261 325
rect 264 323 266 325
rect 269 323 271 325
rect 274 323 276 325
rect 279 323 281 325
rect 284 323 286 325
rect 289 323 291 325
rect 294 323 296 325
rect 4 313 6 315
rect 9 313 11 315
rect 14 313 16 315
rect 19 313 21 315
rect 24 313 26 315
rect 29 313 31 315
rect 34 313 36 315
rect 39 313 41 315
rect 44 313 46 315
rect 49 313 51 315
rect 54 313 56 315
rect 59 313 61 315
rect 64 313 66 315
rect 69 313 71 315
rect 74 313 76 315
rect 79 313 81 315
rect 84 313 86 315
rect 89 313 91 315
rect 94 313 96 315
rect 99 313 101 315
rect 104 313 106 315
rect 109 313 111 315
rect 114 313 116 315
rect 119 313 121 315
rect 124 313 126 315
rect 129 313 131 315
rect 134 313 136 315
rect 139 313 141 315
rect 144 313 146 315
rect 149 313 151 315
rect 154 313 156 315
rect 159 313 161 315
rect 164 313 166 315
rect 169 313 171 315
rect 174 313 176 315
rect 179 313 181 315
rect 184 313 186 315
rect 189 313 191 315
rect 194 313 196 315
rect 199 313 201 315
rect 204 313 206 315
rect 209 313 211 315
rect 214 313 216 315
rect 219 313 221 315
rect 224 313 226 315
rect 229 313 231 315
rect 234 313 236 315
rect 239 313 241 315
rect 244 313 246 315
rect 249 313 251 315
rect 254 313 256 315
rect 259 313 261 315
rect 264 313 266 315
rect 269 313 271 315
rect 274 313 276 315
rect 279 313 281 315
rect 284 313 286 315
rect 289 313 291 315
rect 294 313 296 315
rect 4 303 6 305
rect 9 303 11 305
rect 14 303 16 305
rect 19 303 21 305
rect 24 303 26 305
rect 29 303 31 305
rect 34 303 36 305
rect 39 303 41 305
rect 44 303 46 305
rect 49 303 51 305
rect 54 303 56 305
rect 59 303 61 305
rect 64 303 66 305
rect 69 303 71 305
rect 74 303 76 305
rect 79 303 81 305
rect 84 303 86 305
rect 89 303 91 305
rect 94 303 96 305
rect 99 303 101 305
rect 104 303 106 305
rect 109 303 111 305
rect 114 303 116 305
rect 119 303 121 305
rect 124 303 126 305
rect 129 303 131 305
rect 134 303 136 305
rect 139 303 141 305
rect 144 303 146 305
rect 149 303 151 305
rect 154 303 156 305
rect 159 303 161 305
rect 164 303 166 305
rect 169 303 171 305
rect 174 303 176 305
rect 179 303 181 305
rect 184 303 186 305
rect 189 303 191 305
rect 194 303 196 305
rect 199 303 201 305
rect 204 303 206 305
rect 209 303 211 305
rect 214 303 216 305
rect 219 303 221 305
rect 224 303 226 305
rect 229 303 231 305
rect 234 303 236 305
rect 239 303 241 305
rect 244 303 246 305
rect 249 303 251 305
rect 254 303 256 305
rect 259 303 261 305
rect 264 303 266 305
rect 269 303 271 305
rect 274 303 276 305
rect 279 303 281 305
rect 284 303 286 305
rect 289 303 291 305
rect 294 303 296 305
rect 4 293 6 295
rect 9 293 11 295
rect 14 293 16 295
rect 19 293 21 295
rect 24 293 26 295
rect 29 293 31 295
rect 34 293 36 295
rect 39 293 41 295
rect 44 293 46 295
rect 49 293 51 295
rect 54 293 56 295
rect 59 293 61 295
rect 64 293 66 295
rect 69 293 71 295
rect 74 293 76 295
rect 79 293 81 295
rect 84 293 86 295
rect 89 293 91 295
rect 94 293 96 295
rect 99 293 101 295
rect 104 293 106 295
rect 109 293 111 295
rect 114 293 116 295
rect 119 293 121 295
rect 124 293 126 295
rect 129 293 131 295
rect 134 293 136 295
rect 139 293 141 295
rect 144 293 146 295
rect 149 293 151 295
rect 154 293 156 295
rect 159 293 161 295
rect 164 293 166 295
rect 169 293 171 295
rect 174 293 176 295
rect 179 293 181 295
rect 184 293 186 295
rect 189 293 191 295
rect 194 293 196 295
rect 199 293 201 295
rect 204 293 206 295
rect 209 293 211 295
rect 214 293 216 295
rect 219 293 221 295
rect 224 293 226 295
rect 229 293 231 295
rect 234 293 236 295
rect 239 293 241 295
rect 244 293 246 295
rect 249 293 251 295
rect 254 293 256 295
rect 259 293 261 295
rect 264 293 266 295
rect 269 293 271 295
rect 274 293 276 295
rect 279 293 281 295
rect 284 293 286 295
rect 289 293 291 295
rect 294 293 296 295
rect 4 283 6 285
rect 9 283 11 285
rect 14 283 16 285
rect 19 283 21 285
rect 24 283 26 285
rect 29 283 31 285
rect 34 283 36 285
rect 39 283 41 285
rect 44 283 46 285
rect 49 283 51 285
rect 54 283 56 285
rect 59 283 61 285
rect 64 283 66 285
rect 69 283 71 285
rect 74 283 76 285
rect 79 283 81 285
rect 84 283 86 285
rect 89 283 91 285
rect 94 283 96 285
rect 99 283 101 285
rect 104 283 106 285
rect 109 283 111 285
rect 114 283 116 285
rect 119 283 121 285
rect 124 283 126 285
rect 129 283 131 285
rect 134 283 136 285
rect 139 283 141 285
rect 144 283 146 285
rect 149 283 151 285
rect 154 283 156 285
rect 159 283 161 285
rect 164 283 166 285
rect 169 283 171 285
rect 174 283 176 285
rect 179 283 181 285
rect 184 283 186 285
rect 189 283 191 285
rect 194 283 196 285
rect 199 283 201 285
rect 204 283 206 285
rect 209 283 211 285
rect 214 283 216 285
rect 219 283 221 285
rect 224 283 226 285
rect 229 283 231 285
rect 234 283 236 285
rect 239 283 241 285
rect 244 283 246 285
rect 249 283 251 285
rect 254 283 256 285
rect 259 283 261 285
rect 264 283 266 285
rect 269 283 271 285
rect 274 283 276 285
rect 279 283 281 285
rect 284 283 286 285
rect 289 283 291 285
rect 294 283 296 285
rect 4 273 6 275
rect 9 273 11 275
rect 14 273 16 275
rect 19 273 21 275
rect 24 273 26 275
rect 29 273 31 275
rect 34 273 36 275
rect 39 273 41 275
rect 44 273 46 275
rect 49 273 51 275
rect 54 273 56 275
rect 59 273 61 275
rect 64 273 66 275
rect 69 273 71 275
rect 74 273 76 275
rect 79 273 81 275
rect 84 273 86 275
rect 89 273 91 275
rect 94 273 96 275
rect 99 273 101 275
rect 104 273 106 275
rect 109 273 111 275
rect 114 273 116 275
rect 119 273 121 275
rect 124 273 126 275
rect 129 273 131 275
rect 134 273 136 275
rect 139 273 141 275
rect 144 273 146 275
rect 149 273 151 275
rect 154 273 156 275
rect 159 273 161 275
rect 164 273 166 275
rect 169 273 171 275
rect 174 273 176 275
rect 179 273 181 275
rect 184 273 186 275
rect 189 273 191 275
rect 194 273 196 275
rect 199 273 201 275
rect 204 273 206 275
rect 209 273 211 275
rect 214 273 216 275
rect 219 273 221 275
rect 224 273 226 275
rect 229 273 231 275
rect 234 273 236 275
rect 239 273 241 275
rect 244 273 246 275
rect 249 273 251 275
rect 254 273 256 275
rect 259 273 261 275
rect 264 273 266 275
rect 269 273 271 275
rect 274 273 276 275
rect 279 273 281 275
rect 284 273 286 275
rect 289 273 291 275
rect 294 273 296 275
rect 4 263 6 265
rect 9 263 11 265
rect 14 263 16 265
rect 19 263 21 265
rect 24 263 26 265
rect 29 263 31 265
rect 34 263 36 265
rect 39 263 41 265
rect 44 263 46 265
rect 49 263 51 265
rect 54 263 56 265
rect 59 263 61 265
rect 64 263 66 265
rect 69 263 71 265
rect 74 263 76 265
rect 79 263 81 265
rect 84 263 86 265
rect 89 263 91 265
rect 94 263 96 265
rect 99 263 101 265
rect 104 263 106 265
rect 109 263 111 265
rect 114 263 116 265
rect 119 263 121 265
rect 124 263 126 265
rect 129 263 131 265
rect 134 263 136 265
rect 139 263 141 265
rect 144 263 146 265
rect 149 263 151 265
rect 154 263 156 265
rect 159 263 161 265
rect 164 263 166 265
rect 169 263 171 265
rect 174 263 176 265
rect 179 263 181 265
rect 184 263 186 265
rect 189 263 191 265
rect 194 263 196 265
rect 199 263 201 265
rect 204 263 206 265
rect 209 263 211 265
rect 214 263 216 265
rect 219 263 221 265
rect 224 263 226 265
rect 229 263 231 265
rect 234 263 236 265
rect 239 263 241 265
rect 244 263 246 265
rect 249 263 251 265
rect 254 263 256 265
rect 259 263 261 265
rect 264 263 266 265
rect 269 263 271 265
rect 274 263 276 265
rect 279 263 281 265
rect 284 263 286 265
rect 289 263 291 265
rect 294 263 296 265
rect 3 253 5 255
rect 9 253 11 255
rect 14 253 16 255
rect 19 253 21 255
rect 24 253 26 255
rect 29 253 31 255
rect 34 253 36 255
rect 39 253 41 255
rect 44 253 46 255
rect 49 253 51 255
rect 54 253 56 255
rect 59 253 61 255
rect 64 253 66 255
rect 69 253 71 255
rect 74 253 76 255
rect 79 253 81 255
rect 84 253 86 255
rect 89 253 91 255
rect 94 253 96 255
rect 99 253 101 255
rect 104 253 106 255
rect 109 253 111 255
rect 114 253 116 255
rect 119 253 121 255
rect 124 253 126 255
rect 129 253 131 255
rect 134 253 136 255
rect 139 253 141 255
rect 144 253 146 255
rect 149 253 151 255
rect 154 253 156 255
rect 159 253 161 255
rect 164 253 166 255
rect 169 253 171 255
rect 174 253 176 255
rect 179 253 181 255
rect 184 253 186 255
rect 189 253 191 255
rect 194 253 196 255
rect 199 253 201 255
rect 204 253 206 255
rect 209 253 211 255
rect 214 253 216 255
rect 219 253 221 255
rect 224 253 226 255
rect 229 253 231 255
rect 234 253 236 255
rect 239 253 241 255
rect 244 253 246 255
rect 249 253 251 255
rect 254 253 256 255
rect 259 253 261 255
rect 264 253 266 255
rect 269 253 271 255
rect 274 253 276 255
rect 279 253 281 255
rect 284 253 286 255
rect 289 253 291 255
rect 295 253 297 255
rect 3 248 5 250
rect 295 248 297 250
rect 3 243 5 245
rect 295 243 297 245
rect 203 240 205 242
rect 208 240 210 242
rect 213 240 215 242
rect 218 240 220 242
rect 223 240 225 242
rect 228 240 230 242
rect 233 240 235 242
rect 238 240 240 242
rect 243 240 245 242
rect 248 240 250 242
rect 253 240 255 242
rect 258 240 260 242
rect 263 240 265 242
rect 268 240 270 242
rect 273 240 275 242
rect 278 240 280 242
rect 3 238 5 240
rect 20 237 22 239
rect 25 237 27 239
rect 30 237 32 239
rect 35 237 37 239
rect 40 237 42 239
rect 45 237 47 239
rect 50 237 52 239
rect 55 237 57 239
rect 60 237 62 239
rect 65 237 67 239
rect 70 237 72 239
rect 75 237 77 239
rect 80 237 82 239
rect 85 237 87 239
rect 90 237 92 239
rect 95 237 97 239
rect 295 238 297 240
rect 203 235 205 237
rect 208 235 210 237
rect 213 235 215 237
rect 218 235 220 237
rect 223 235 225 237
rect 228 235 230 237
rect 233 235 235 237
rect 238 235 240 237
rect 243 235 245 237
rect 248 235 250 237
rect 253 235 255 237
rect 258 235 260 237
rect 263 235 265 237
rect 268 235 270 237
rect 273 235 275 237
rect 278 235 280 237
rect 3 233 5 235
rect 295 233 297 235
rect 3 228 5 230
rect 25 229 27 231
rect 40 229 42 231
rect 45 229 47 231
rect 50 229 52 231
rect 55 229 57 231
rect 60 229 62 231
rect 65 229 67 231
rect 70 229 72 231
rect 75 229 77 231
rect 80 229 82 231
rect 85 229 87 231
rect 90 229 92 231
rect 95 229 97 231
rect 203 229 205 231
rect 208 229 210 231
rect 213 229 215 231
rect 218 229 220 231
rect 223 229 225 231
rect 228 229 230 231
rect 233 229 235 231
rect 238 229 240 231
rect 243 229 245 231
rect 248 229 250 231
rect 253 229 255 231
rect 258 229 260 231
rect 278 229 280 231
rect 295 228 297 230
rect 3 223 5 225
rect 25 224 27 226
rect 42 223 44 225
rect 47 223 49 225
rect 52 223 54 225
rect 57 223 59 225
rect 62 223 64 225
rect 67 223 69 225
rect 72 223 74 225
rect 77 223 79 225
rect 82 223 84 225
rect 87 223 89 225
rect 92 223 94 225
rect 206 223 208 225
rect 211 223 213 225
rect 216 223 218 225
rect 221 223 223 225
rect 226 223 228 225
rect 231 223 233 225
rect 236 223 238 225
rect 241 223 243 225
rect 246 223 248 225
rect 251 223 253 225
rect 256 223 258 225
rect 278 224 280 226
rect 295 223 297 225
rect 3 218 5 220
rect 25 219 27 221
rect 146 219 148 221
rect 151 219 153 221
rect 278 219 280 221
rect 295 218 297 220
rect 3 213 5 215
rect 25 214 27 216
rect 33 213 35 215
rect 265 213 267 215
rect 278 214 280 216
rect 295 213 297 215
rect 146 211 148 213
rect 151 211 153 213
rect 3 208 5 210
rect 25 209 27 211
rect 33 208 35 210
rect 265 208 267 210
rect 278 209 280 211
rect 295 208 297 210
rect 3 203 5 205
rect 25 204 27 206
rect 33 203 35 205
rect 146 203 148 205
rect 151 203 153 205
rect 265 203 267 205
rect 278 204 280 206
rect 295 203 297 205
rect 3 198 5 200
rect 25 199 27 201
rect 33 198 35 200
rect 265 198 267 200
rect 278 199 280 201
rect 295 198 297 200
rect 57 196 59 198
rect 62 196 64 198
rect 67 196 69 198
rect 72 196 74 198
rect 77 196 79 198
rect 82 196 84 198
rect 87 196 89 198
rect 92 196 94 198
rect 97 196 99 198
rect 102 196 104 198
rect 107 196 109 198
rect 112 196 114 198
rect 117 196 119 198
rect 181 196 183 198
rect 186 196 188 198
rect 191 196 193 198
rect 196 196 198 198
rect 201 196 203 198
rect 206 196 208 198
rect 211 196 213 198
rect 216 196 218 198
rect 221 196 223 198
rect 226 196 228 198
rect 231 196 233 198
rect 236 196 238 198
rect 241 196 243 198
rect 3 193 5 195
rect 25 194 27 196
rect 33 193 35 195
rect 265 193 267 195
rect 278 194 280 196
rect 295 193 297 195
rect 3 188 5 190
rect 25 189 27 191
rect 57 190 59 192
rect 62 190 64 192
rect 67 190 69 192
rect 72 190 74 192
rect 77 190 79 192
rect 82 190 84 192
rect 87 190 89 192
rect 92 190 94 192
rect 97 190 99 192
rect 102 190 104 192
rect 107 190 109 192
rect 112 190 114 192
rect 117 190 119 192
rect 181 190 183 192
rect 186 190 188 192
rect 191 190 193 192
rect 196 190 198 192
rect 201 190 203 192
rect 206 190 208 192
rect 211 190 213 192
rect 216 190 218 192
rect 221 190 223 192
rect 226 190 228 192
rect 231 190 233 192
rect 236 190 238 192
rect 241 190 243 192
rect 33 188 35 190
rect 265 188 267 190
rect 278 189 280 191
rect 295 188 297 190
rect 3 183 5 185
rect 25 184 27 186
rect 33 183 35 185
rect 265 183 267 185
rect 278 184 280 186
rect 295 183 297 185
rect 3 178 5 180
rect 25 179 27 181
rect 33 178 35 180
rect 265 178 267 180
rect 278 179 280 181
rect 295 178 297 180
rect 3 173 5 175
rect 25 174 27 176
rect 33 173 35 175
rect 265 173 267 175
rect 278 174 280 176
rect 295 173 297 175
rect 3 168 5 170
rect 25 169 27 171
rect 33 168 35 170
rect 265 168 267 170
rect 278 169 280 171
rect 295 168 297 170
rect 3 163 5 165
rect 25 164 27 166
rect 33 163 35 165
rect 42 163 44 165
rect 47 163 49 165
rect 52 163 54 165
rect 57 163 59 165
rect 62 163 64 165
rect 67 163 69 165
rect 72 163 74 165
rect 77 163 79 165
rect 82 163 84 165
rect 87 163 89 165
rect 92 163 94 165
rect 97 163 99 165
rect 102 163 104 165
rect 107 163 109 165
rect 112 163 114 165
rect 117 163 119 165
rect 181 163 183 165
rect 186 163 188 165
rect 191 163 193 165
rect 196 163 198 165
rect 201 163 203 165
rect 206 163 208 165
rect 211 163 213 165
rect 216 163 218 165
rect 221 163 223 165
rect 226 163 228 165
rect 231 163 233 165
rect 236 163 238 165
rect 241 163 243 165
rect 246 163 248 165
rect 251 163 253 165
rect 256 163 258 165
rect 265 163 267 165
rect 278 164 280 166
rect 295 163 297 165
rect 3 158 5 160
rect 25 159 27 161
rect 33 158 35 160
rect 42 157 44 159
rect 47 157 49 159
rect 52 157 54 159
rect 57 157 59 159
rect 62 157 64 159
rect 67 157 69 159
rect 72 157 74 159
rect 77 157 79 159
rect 82 157 84 159
rect 87 157 89 159
rect 92 157 94 159
rect 97 157 99 159
rect 102 157 104 159
rect 107 157 109 159
rect 112 157 114 159
rect 117 157 119 159
rect 181 157 183 159
rect 186 157 188 159
rect 191 157 193 159
rect 196 157 198 159
rect 201 157 203 159
rect 206 157 208 159
rect 211 157 213 159
rect 216 157 218 159
rect 221 157 223 159
rect 226 157 228 159
rect 231 157 233 159
rect 236 157 238 159
rect 241 157 243 159
rect 246 157 248 159
rect 251 157 253 159
rect 256 157 258 159
rect 265 158 267 160
rect 278 159 280 161
rect 295 158 297 160
rect 3 153 5 155
rect 25 154 27 156
rect 33 153 35 155
rect 265 153 267 155
rect 278 154 280 156
rect 295 153 297 155
rect 3 148 5 150
rect 25 149 27 151
rect 33 148 35 150
rect 265 148 267 150
rect 278 149 280 151
rect 295 148 297 150
rect 3 143 5 145
rect 25 144 27 146
rect 33 143 35 145
rect 265 143 267 145
rect 278 144 280 146
rect 295 143 297 145
rect 3 138 5 140
rect 25 139 27 141
rect 33 138 35 140
rect 265 138 267 140
rect 278 139 280 141
rect 295 138 297 140
rect 3 133 5 135
rect 25 134 27 136
rect 33 133 35 135
rect 265 133 267 135
rect 278 134 280 136
rect 295 133 297 135
rect 3 128 5 130
rect 25 129 27 131
rect 57 130 59 132
rect 62 130 64 132
rect 67 130 69 132
rect 72 130 74 132
rect 77 130 79 132
rect 82 130 84 132
rect 87 130 89 132
rect 92 130 94 132
rect 97 130 99 132
rect 102 130 104 132
rect 107 130 109 132
rect 112 130 114 132
rect 117 130 119 132
rect 146 131 148 133
rect 151 131 153 133
rect 181 130 183 132
rect 186 130 188 132
rect 191 130 193 132
rect 196 130 198 132
rect 201 130 203 132
rect 206 130 208 132
rect 211 130 213 132
rect 216 130 218 132
rect 221 130 223 132
rect 226 130 228 132
rect 231 130 233 132
rect 236 130 238 132
rect 241 130 243 132
rect 33 128 35 130
rect 265 128 267 130
rect 278 129 280 131
rect 295 128 297 130
rect 3 123 5 125
rect 25 124 27 126
rect 57 125 59 127
rect 62 125 64 127
rect 67 125 69 127
rect 72 125 74 127
rect 77 125 79 127
rect 82 125 84 127
rect 87 125 89 127
rect 92 125 94 127
rect 97 125 99 127
rect 102 125 104 127
rect 107 125 109 127
rect 112 125 114 127
rect 117 125 119 127
rect 181 125 183 127
rect 186 125 188 127
rect 191 125 193 127
rect 196 125 198 127
rect 201 125 203 127
rect 206 125 208 127
rect 211 125 213 127
rect 216 125 218 127
rect 221 125 223 127
rect 226 125 228 127
rect 231 125 233 127
rect 236 125 238 127
rect 241 125 243 127
rect 33 123 35 125
rect 146 123 148 125
rect 151 123 153 125
rect 265 123 267 125
rect 278 124 280 126
rect 295 123 297 125
rect 3 118 5 120
rect 25 119 27 121
rect 33 118 35 120
rect 265 118 267 120
rect 278 119 280 121
rect 295 118 297 120
rect 3 113 5 115
rect 25 114 27 116
rect 33 113 35 115
rect 265 113 267 115
rect 278 114 280 116
rect 295 113 297 115
rect 3 108 5 110
rect 25 109 27 111
rect 33 108 35 110
rect 265 108 267 110
rect 278 109 280 111
rect 295 108 297 110
rect 3 103 5 105
rect 25 104 27 106
rect 33 103 35 105
rect 265 103 267 105
rect 278 104 280 106
rect 295 103 297 105
rect 3 98 5 100
rect 25 99 27 101
rect 33 98 35 100
rect 42 98 44 100
rect 47 98 49 100
rect 52 98 54 100
rect 57 98 59 100
rect 62 98 64 100
rect 67 98 69 100
rect 72 98 74 100
rect 77 98 79 100
rect 82 98 84 100
rect 87 98 89 100
rect 92 98 94 100
rect 97 98 99 100
rect 102 98 104 100
rect 107 98 109 100
rect 112 98 114 100
rect 117 98 119 100
rect 181 98 183 100
rect 186 98 188 100
rect 191 98 193 100
rect 196 98 198 100
rect 201 98 203 100
rect 206 98 208 100
rect 211 98 213 100
rect 216 98 218 100
rect 221 98 223 100
rect 226 98 228 100
rect 231 98 233 100
rect 236 98 238 100
rect 241 98 243 100
rect 246 98 248 100
rect 251 98 253 100
rect 256 98 258 100
rect 265 98 267 100
rect 278 99 280 101
rect 295 98 297 100
rect 3 93 5 95
rect 25 94 27 96
rect 33 93 35 95
rect 42 92 44 94
rect 47 92 49 94
rect 52 92 54 94
rect 57 92 59 94
rect 62 92 64 94
rect 67 92 69 94
rect 72 92 74 94
rect 77 92 79 94
rect 82 92 84 94
rect 87 92 89 94
rect 92 92 94 94
rect 97 92 99 94
rect 102 92 104 94
rect 107 92 109 94
rect 112 92 114 94
rect 117 92 119 94
rect 181 92 183 94
rect 186 92 188 94
rect 191 92 193 94
rect 196 92 198 94
rect 201 92 203 94
rect 206 92 208 94
rect 211 92 213 94
rect 216 92 218 94
rect 221 92 223 94
rect 226 92 228 94
rect 231 92 233 94
rect 236 92 238 94
rect 241 92 243 94
rect 246 92 248 94
rect 251 92 253 94
rect 256 92 258 94
rect 265 93 267 95
rect 278 94 280 96
rect 295 93 297 95
rect 3 88 5 90
rect 25 89 27 91
rect 33 88 35 90
rect 265 88 267 90
rect 278 89 280 91
rect 295 88 297 90
rect 3 83 5 85
rect 25 84 27 86
rect 33 83 35 85
rect 265 83 267 85
rect 278 84 280 86
rect 295 83 297 85
rect 3 78 5 80
rect 25 79 27 81
rect 33 78 35 80
rect 265 78 267 80
rect 278 79 280 81
rect 295 78 297 80
rect 3 73 5 75
rect 25 74 27 76
rect 33 73 35 75
rect 265 73 267 75
rect 278 74 280 76
rect 295 73 297 75
rect 3 68 5 70
rect 25 69 27 71
rect 33 68 35 70
rect 265 68 267 70
rect 278 69 280 71
rect 295 68 297 70
rect 3 63 5 65
rect 25 64 27 66
rect 57 65 59 67
rect 62 65 64 67
rect 67 65 69 67
rect 72 65 74 67
rect 77 65 79 67
rect 82 65 84 67
rect 87 65 89 67
rect 92 65 94 67
rect 97 65 99 67
rect 102 65 104 67
rect 107 65 109 67
rect 112 65 114 67
rect 117 65 119 67
rect 181 65 183 67
rect 186 65 188 67
rect 191 65 193 67
rect 196 65 198 67
rect 201 65 203 67
rect 206 65 208 67
rect 211 65 213 67
rect 216 65 218 67
rect 221 65 223 67
rect 226 65 228 67
rect 231 65 233 67
rect 236 65 238 67
rect 241 65 243 67
rect 33 63 35 65
rect 265 63 267 65
rect 278 64 280 66
rect 295 63 297 65
rect 3 58 5 60
rect 25 59 27 61
rect 57 60 59 62
rect 62 60 64 62
rect 67 60 69 62
rect 72 60 74 62
rect 77 60 79 62
rect 82 60 84 62
rect 87 60 89 62
rect 92 60 94 62
rect 97 60 99 62
rect 102 60 104 62
rect 107 60 109 62
rect 112 60 114 62
rect 117 60 119 62
rect 33 58 35 60
rect 146 59 148 61
rect 151 59 153 61
rect 181 60 183 62
rect 186 60 188 62
rect 191 60 193 62
rect 196 60 198 62
rect 201 60 203 62
rect 206 60 208 62
rect 211 60 213 62
rect 216 60 218 62
rect 221 60 223 62
rect 226 60 228 62
rect 231 60 233 62
rect 236 60 238 62
rect 241 60 243 62
rect 265 58 267 60
rect 278 59 280 61
rect 295 58 297 60
rect 3 53 5 55
rect 25 54 27 56
rect 33 53 35 55
rect 265 53 267 55
rect 278 54 280 56
rect 295 53 297 55
rect 146 51 148 53
rect 151 51 153 53
rect 3 48 5 50
rect 25 49 27 51
rect 33 48 35 50
rect 265 48 267 50
rect 278 49 280 51
rect 295 48 297 50
rect 3 43 5 45
rect 25 44 27 46
rect 33 43 35 45
rect 146 43 148 45
rect 151 43 153 45
rect 265 43 267 45
rect 278 44 280 46
rect 295 43 297 45
rect 3 38 5 40
rect 25 39 27 41
rect 278 39 280 41
rect 295 38 297 40
rect 3 33 5 35
rect 25 34 27 36
rect 146 35 148 37
rect 151 35 153 37
rect 42 33 44 35
rect 47 33 49 35
rect 52 33 54 35
rect 57 33 59 35
rect 62 33 64 35
rect 67 33 69 35
rect 72 33 74 35
rect 77 33 79 35
rect 82 33 84 35
rect 87 33 89 35
rect 92 33 94 35
rect 206 33 208 35
rect 211 33 213 35
rect 216 33 218 35
rect 221 33 223 35
rect 226 33 228 35
rect 231 33 233 35
rect 236 33 238 35
rect 241 33 243 35
rect 246 33 248 35
rect 251 33 253 35
rect 256 33 258 35
rect 278 34 280 36
rect 295 33 297 35
rect 3 28 5 30
rect 25 29 27 31
rect 278 29 280 31
rect 295 28 297 30
rect 3 23 5 25
rect 20 23 22 25
rect 25 23 27 25
rect 30 23 32 25
rect 35 23 37 25
rect 40 23 42 25
rect 45 23 47 25
rect 50 23 52 25
rect 55 23 57 25
rect 60 23 62 25
rect 65 23 67 25
rect 70 23 72 25
rect 75 23 77 25
rect 80 23 82 25
rect 85 23 87 25
rect 90 23 92 25
rect 95 23 97 25
rect 203 23 205 25
rect 208 23 210 25
rect 213 23 215 25
rect 218 23 220 25
rect 223 23 225 25
rect 228 23 230 25
rect 233 23 235 25
rect 238 23 240 25
rect 243 23 245 25
rect 248 23 250 25
rect 253 23 255 25
rect 258 23 260 25
rect 263 23 265 25
rect 268 23 270 25
rect 273 23 275 25
rect 278 23 280 25
rect 295 23 297 25
rect 3 18 5 20
rect 295 18 297 20
rect 3 13 5 15
rect 295 13 297 15
rect 3 8 5 10
rect 295 8 297 10
rect 3 3 5 5
rect 9 3 11 5
rect 14 3 16 5
rect 19 3 21 5
rect 24 3 26 5
rect 29 3 31 5
rect 34 3 36 5
rect 39 3 41 5
rect 44 3 46 5
rect 49 3 51 5
rect 54 3 56 5
rect 59 3 61 5
rect 64 3 66 5
rect 69 3 71 5
rect 74 3 76 5
rect 79 3 81 5
rect 84 3 86 5
rect 89 3 91 5
rect 204 3 206 5
rect 209 3 211 5
rect 214 3 216 5
rect 219 3 221 5
rect 224 3 226 5
rect 229 3 231 5
rect 234 3 236 5
rect 239 3 241 5
rect 244 3 246 5
rect 249 3 251 5
rect 254 3 256 5
rect 259 3 261 5
rect 264 3 266 5
rect 269 3 271 5
rect 274 3 276 5
rect 279 3 281 5
rect 284 3 286 5
rect 289 3 291 5
rect 295 3 297 5
<< metal1 >>
rect 20 740 280 1000
rect 62 730 238 740
rect 72 720 228 730
rect 82 710 218 720
rect 92 700 208 710
rect 0 659 99 670
rect 0 419 10 659
rect 102 650 198 700
rect 201 659 300 670
rect 50 649 280 650
rect 21 433 280 649
rect 102 424 198 433
rect 0 344 99 419
rect 102 340 140 424
rect 143 344 157 421
rect 160 340 198 424
rect 289 419 300 659
rect 201 344 300 419
rect 102 326 198 340
rect 0 251 300 326
rect 0 7 8 251
rect 14 210 99 245
rect 102 229 198 251
rect 14 178 53 210
rect 102 207 142 229
rect 56 199 142 207
rect 145 202 154 226
rect 157 207 198 229
rect 201 210 286 245
rect 157 199 244 207
rect 56 181 244 199
rect 14 144 120 178
rect 14 113 53 144
rect 123 141 177 181
rect 247 178 286 210
rect 180 144 286 178
rect 56 137 244 141
rect 56 119 142 137
rect 145 122 154 134
rect 157 119 244 137
rect 56 116 244 119
rect 14 79 120 113
rect 14 48 53 79
rect 123 76 177 116
rect 247 113 286 144
rect 180 79 286 113
rect 56 69 244 76
rect 56 51 142 69
rect 14 13 99 48
rect 102 27 142 51
rect 145 30 154 66
rect 157 51 244 69
rect 157 27 198 51
rect 247 48 286 79
rect 0 -1 99 7
rect 102 -12 198 27
rect 201 13 286 48
rect 292 7 300 251
rect 201 -1 300 7
<< metal2 >>
rect 20 740 280 1000
rect 0 440 300 670
rect 0 344 300 424
rect 0 246 300 326
rect 0 6 300 229
rect 0 -1 98 6
rect 202 -1 300 6
<< gv1 >>
rect 41 977 43 979
rect 53 977 55 979
rect 65 977 67 979
rect 77 977 79 979
rect 89 977 91 979
rect 101 977 103 979
rect 113 977 115 979
rect 125 977 127 979
rect 137 977 139 979
rect 149 977 151 979
rect 161 977 163 979
rect 173 977 175 979
rect 185 977 187 979
rect 197 977 199 979
rect 209 977 211 979
rect 221 977 223 979
rect 233 977 235 979
rect 245 977 247 979
rect 257 977 259 979
rect 41 965 43 967
rect 53 965 55 967
rect 65 965 67 967
rect 77 965 79 967
rect 89 965 91 967
rect 101 965 103 967
rect 113 965 115 967
rect 125 965 127 967
rect 137 965 139 967
rect 149 965 151 967
rect 161 965 163 967
rect 173 965 175 967
rect 185 965 187 967
rect 197 965 199 967
rect 209 965 211 967
rect 221 965 223 967
rect 233 965 235 967
rect 245 965 247 967
rect 257 965 259 967
rect 41 953 43 955
rect 53 953 55 955
rect 65 953 67 955
rect 77 953 79 955
rect 89 953 91 955
rect 101 953 103 955
rect 113 953 115 955
rect 125 953 127 955
rect 137 953 139 955
rect 149 953 151 955
rect 161 953 163 955
rect 173 953 175 955
rect 185 953 187 955
rect 197 953 199 955
rect 209 953 211 955
rect 221 953 223 955
rect 233 953 235 955
rect 245 953 247 955
rect 257 953 259 955
rect 41 941 43 943
rect 53 941 55 943
rect 65 941 67 943
rect 77 941 79 943
rect 89 941 91 943
rect 101 941 103 943
rect 113 941 115 943
rect 125 941 127 943
rect 137 941 139 943
rect 149 941 151 943
rect 161 941 163 943
rect 173 941 175 943
rect 185 941 187 943
rect 197 941 199 943
rect 209 941 211 943
rect 221 941 223 943
rect 233 941 235 943
rect 245 941 247 943
rect 257 941 259 943
rect 41 929 43 931
rect 53 929 55 931
rect 65 929 67 931
rect 77 929 79 931
rect 89 929 91 931
rect 101 929 103 931
rect 113 929 115 931
rect 125 929 127 931
rect 137 929 139 931
rect 149 929 151 931
rect 161 929 163 931
rect 173 929 175 931
rect 185 929 187 931
rect 197 929 199 931
rect 209 929 211 931
rect 221 929 223 931
rect 233 929 235 931
rect 245 929 247 931
rect 257 929 259 931
rect 41 917 43 919
rect 53 917 55 919
rect 65 917 67 919
rect 77 917 79 919
rect 89 917 91 919
rect 101 917 103 919
rect 113 917 115 919
rect 125 917 127 919
rect 137 917 139 919
rect 149 917 151 919
rect 161 917 163 919
rect 173 917 175 919
rect 185 917 187 919
rect 197 917 199 919
rect 209 917 211 919
rect 221 917 223 919
rect 233 917 235 919
rect 245 917 247 919
rect 257 917 259 919
rect 41 905 43 907
rect 53 905 55 907
rect 65 905 67 907
rect 77 905 79 907
rect 89 905 91 907
rect 101 905 103 907
rect 113 905 115 907
rect 125 905 127 907
rect 137 905 139 907
rect 149 905 151 907
rect 161 905 163 907
rect 173 905 175 907
rect 185 905 187 907
rect 197 905 199 907
rect 209 905 211 907
rect 221 905 223 907
rect 233 905 235 907
rect 245 905 247 907
rect 257 905 259 907
rect 41 893 43 895
rect 53 893 55 895
rect 65 893 67 895
rect 77 893 79 895
rect 89 893 91 895
rect 101 893 103 895
rect 113 893 115 895
rect 125 893 127 895
rect 137 893 139 895
rect 149 893 151 895
rect 161 893 163 895
rect 173 893 175 895
rect 185 893 187 895
rect 197 893 199 895
rect 209 893 211 895
rect 221 893 223 895
rect 233 893 235 895
rect 245 893 247 895
rect 257 893 259 895
rect 41 881 43 883
rect 53 881 55 883
rect 65 881 67 883
rect 77 881 79 883
rect 89 881 91 883
rect 101 881 103 883
rect 113 881 115 883
rect 125 881 127 883
rect 137 881 139 883
rect 149 881 151 883
rect 161 881 163 883
rect 173 881 175 883
rect 185 881 187 883
rect 197 881 199 883
rect 209 881 211 883
rect 221 881 223 883
rect 233 881 235 883
rect 245 881 247 883
rect 257 881 259 883
rect 41 869 43 871
rect 53 869 55 871
rect 65 869 67 871
rect 77 869 79 871
rect 89 869 91 871
rect 101 869 103 871
rect 113 869 115 871
rect 125 869 127 871
rect 137 869 139 871
rect 149 869 151 871
rect 161 869 163 871
rect 173 869 175 871
rect 185 869 187 871
rect 197 869 199 871
rect 209 869 211 871
rect 221 869 223 871
rect 233 869 235 871
rect 245 869 247 871
rect 257 869 259 871
rect 41 857 43 859
rect 53 857 55 859
rect 65 857 67 859
rect 77 857 79 859
rect 89 857 91 859
rect 101 857 103 859
rect 113 857 115 859
rect 125 857 127 859
rect 137 857 139 859
rect 149 857 151 859
rect 161 857 163 859
rect 173 857 175 859
rect 185 857 187 859
rect 197 857 199 859
rect 209 857 211 859
rect 221 857 223 859
rect 233 857 235 859
rect 245 857 247 859
rect 257 857 259 859
rect 41 845 43 847
rect 53 845 55 847
rect 65 845 67 847
rect 77 845 79 847
rect 89 845 91 847
rect 101 845 103 847
rect 113 845 115 847
rect 125 845 127 847
rect 137 845 139 847
rect 149 845 151 847
rect 161 845 163 847
rect 173 845 175 847
rect 185 845 187 847
rect 197 845 199 847
rect 209 845 211 847
rect 221 845 223 847
rect 233 845 235 847
rect 245 845 247 847
rect 257 845 259 847
rect 41 833 43 835
rect 53 833 55 835
rect 65 833 67 835
rect 77 833 79 835
rect 89 833 91 835
rect 101 833 103 835
rect 113 833 115 835
rect 125 833 127 835
rect 137 833 139 835
rect 149 833 151 835
rect 161 833 163 835
rect 173 833 175 835
rect 185 833 187 835
rect 197 833 199 835
rect 209 833 211 835
rect 221 833 223 835
rect 233 833 235 835
rect 245 833 247 835
rect 257 833 259 835
rect 41 821 43 823
rect 53 821 55 823
rect 65 821 67 823
rect 77 821 79 823
rect 89 821 91 823
rect 101 821 103 823
rect 113 821 115 823
rect 125 821 127 823
rect 137 821 139 823
rect 149 821 151 823
rect 161 821 163 823
rect 173 821 175 823
rect 185 821 187 823
rect 197 821 199 823
rect 209 821 211 823
rect 221 821 223 823
rect 233 821 235 823
rect 245 821 247 823
rect 257 821 259 823
rect 41 809 43 811
rect 53 809 55 811
rect 65 809 67 811
rect 77 809 79 811
rect 89 809 91 811
rect 101 809 103 811
rect 113 809 115 811
rect 125 809 127 811
rect 137 809 139 811
rect 149 809 151 811
rect 161 809 163 811
rect 173 809 175 811
rect 185 809 187 811
rect 197 809 199 811
rect 209 809 211 811
rect 221 809 223 811
rect 233 809 235 811
rect 245 809 247 811
rect 257 809 259 811
rect 41 797 43 799
rect 53 797 55 799
rect 65 797 67 799
rect 77 797 79 799
rect 89 797 91 799
rect 101 797 103 799
rect 113 797 115 799
rect 125 797 127 799
rect 137 797 139 799
rect 149 797 151 799
rect 161 797 163 799
rect 173 797 175 799
rect 185 797 187 799
rect 197 797 199 799
rect 209 797 211 799
rect 221 797 223 799
rect 233 797 235 799
rect 245 797 247 799
rect 257 797 259 799
rect 41 785 43 787
rect 53 785 55 787
rect 65 785 67 787
rect 77 785 79 787
rect 89 785 91 787
rect 101 785 103 787
rect 113 785 115 787
rect 125 785 127 787
rect 137 785 139 787
rect 149 785 151 787
rect 161 785 163 787
rect 173 785 175 787
rect 185 785 187 787
rect 197 785 199 787
rect 209 785 211 787
rect 221 785 223 787
rect 233 785 235 787
rect 245 785 247 787
rect 257 785 259 787
rect 41 773 43 775
rect 53 773 55 775
rect 65 773 67 775
rect 77 773 79 775
rect 89 773 91 775
rect 101 773 103 775
rect 113 773 115 775
rect 125 773 127 775
rect 137 773 139 775
rect 149 773 151 775
rect 161 773 163 775
rect 173 773 175 775
rect 185 773 187 775
rect 197 773 199 775
rect 209 773 211 775
rect 221 773 223 775
rect 233 773 235 775
rect 245 773 247 775
rect 257 773 259 775
rect 41 761 43 763
rect 53 761 55 763
rect 65 761 67 763
rect 77 761 79 763
rect 89 761 91 763
rect 101 761 103 763
rect 113 761 115 763
rect 125 761 127 763
rect 137 761 139 763
rect 149 761 151 763
rect 161 761 163 763
rect 173 761 175 763
rect 185 761 187 763
rect 197 761 199 763
rect 209 761 211 763
rect 221 761 223 763
rect 233 761 235 763
rect 245 761 247 763
rect 257 761 259 763
rect 24 641 26 643
rect 29 641 31 643
rect 34 641 36 643
rect 39 641 41 643
rect 44 641 46 643
rect 49 641 51 643
rect 54 641 56 643
rect 59 641 61 643
rect 64 641 66 643
rect 69 641 71 643
rect 74 641 76 643
rect 79 641 81 643
rect 84 641 86 643
rect 89 641 91 643
rect 94 641 96 643
rect 99 641 101 643
rect 104 641 106 643
rect 109 641 111 643
rect 114 641 116 643
rect 119 641 121 643
rect 124 641 126 643
rect 129 641 131 643
rect 134 641 136 643
rect 139 641 141 643
rect 144 641 146 643
rect 149 641 151 643
rect 154 641 156 643
rect 159 641 161 643
rect 164 641 166 643
rect 169 641 171 643
rect 174 641 176 643
rect 179 641 181 643
rect 184 641 186 643
rect 189 641 191 643
rect 194 641 196 643
rect 199 641 201 643
rect 204 641 206 643
rect 209 641 211 643
rect 214 641 216 643
rect 219 641 221 643
rect 224 641 226 643
rect 229 641 231 643
rect 234 641 236 643
rect 239 641 241 643
rect 244 641 246 643
rect 249 641 251 643
rect 254 641 256 643
rect 259 641 261 643
rect 264 641 266 643
rect 269 641 271 643
rect 274 641 276 643
rect 24 631 26 633
rect 29 631 31 633
rect 34 631 36 633
rect 39 631 41 633
rect 44 631 46 633
rect 49 631 51 633
rect 54 631 56 633
rect 59 631 61 633
rect 64 631 66 633
rect 69 631 71 633
rect 74 631 76 633
rect 79 631 81 633
rect 84 631 86 633
rect 89 631 91 633
rect 94 631 96 633
rect 99 631 101 633
rect 104 631 106 633
rect 109 631 111 633
rect 114 631 116 633
rect 119 631 121 633
rect 124 631 126 633
rect 129 631 131 633
rect 134 631 136 633
rect 139 631 141 633
rect 144 631 146 633
rect 149 631 151 633
rect 154 631 156 633
rect 159 631 161 633
rect 164 631 166 633
rect 169 631 171 633
rect 174 631 176 633
rect 179 631 181 633
rect 184 631 186 633
rect 189 631 191 633
rect 194 631 196 633
rect 199 631 201 633
rect 204 631 206 633
rect 209 631 211 633
rect 214 631 216 633
rect 219 631 221 633
rect 224 631 226 633
rect 229 631 231 633
rect 234 631 236 633
rect 239 631 241 633
rect 244 631 246 633
rect 249 631 251 633
rect 254 631 256 633
rect 259 631 261 633
rect 264 631 266 633
rect 269 631 271 633
rect 274 631 276 633
rect 24 621 26 623
rect 29 621 31 623
rect 34 621 36 623
rect 39 621 41 623
rect 44 621 46 623
rect 49 621 51 623
rect 54 621 56 623
rect 59 621 61 623
rect 64 621 66 623
rect 69 621 71 623
rect 74 621 76 623
rect 79 621 81 623
rect 84 621 86 623
rect 89 621 91 623
rect 94 621 96 623
rect 99 621 101 623
rect 104 621 106 623
rect 109 621 111 623
rect 114 621 116 623
rect 119 621 121 623
rect 124 621 126 623
rect 129 621 131 623
rect 134 621 136 623
rect 139 621 141 623
rect 144 621 146 623
rect 149 621 151 623
rect 154 621 156 623
rect 159 621 161 623
rect 164 621 166 623
rect 169 621 171 623
rect 174 621 176 623
rect 179 621 181 623
rect 184 621 186 623
rect 189 621 191 623
rect 194 621 196 623
rect 199 621 201 623
rect 204 621 206 623
rect 209 621 211 623
rect 214 621 216 623
rect 219 621 221 623
rect 224 621 226 623
rect 229 621 231 623
rect 234 621 236 623
rect 239 621 241 623
rect 244 621 246 623
rect 249 621 251 623
rect 254 621 256 623
rect 259 621 261 623
rect 264 621 266 623
rect 269 621 271 623
rect 274 621 276 623
rect 24 611 26 613
rect 29 611 31 613
rect 34 611 36 613
rect 39 611 41 613
rect 44 611 46 613
rect 49 611 51 613
rect 54 611 56 613
rect 59 611 61 613
rect 64 611 66 613
rect 69 611 71 613
rect 74 611 76 613
rect 79 611 81 613
rect 84 611 86 613
rect 89 611 91 613
rect 94 611 96 613
rect 99 611 101 613
rect 104 611 106 613
rect 109 611 111 613
rect 114 611 116 613
rect 119 611 121 613
rect 124 611 126 613
rect 129 611 131 613
rect 134 611 136 613
rect 139 611 141 613
rect 144 611 146 613
rect 149 611 151 613
rect 154 611 156 613
rect 159 611 161 613
rect 164 611 166 613
rect 169 611 171 613
rect 174 611 176 613
rect 179 611 181 613
rect 184 611 186 613
rect 189 611 191 613
rect 194 611 196 613
rect 199 611 201 613
rect 204 611 206 613
rect 209 611 211 613
rect 214 611 216 613
rect 219 611 221 613
rect 224 611 226 613
rect 229 611 231 613
rect 234 611 236 613
rect 239 611 241 613
rect 244 611 246 613
rect 249 611 251 613
rect 254 611 256 613
rect 259 611 261 613
rect 264 611 266 613
rect 269 611 271 613
rect 274 611 276 613
rect 24 601 26 603
rect 29 601 31 603
rect 34 601 36 603
rect 39 601 41 603
rect 44 601 46 603
rect 49 601 51 603
rect 54 601 56 603
rect 59 601 61 603
rect 64 601 66 603
rect 69 601 71 603
rect 74 601 76 603
rect 79 601 81 603
rect 84 601 86 603
rect 89 601 91 603
rect 94 601 96 603
rect 99 601 101 603
rect 104 601 106 603
rect 109 601 111 603
rect 114 601 116 603
rect 119 601 121 603
rect 124 601 126 603
rect 129 601 131 603
rect 134 601 136 603
rect 139 601 141 603
rect 144 601 146 603
rect 149 601 151 603
rect 154 601 156 603
rect 159 601 161 603
rect 164 601 166 603
rect 169 601 171 603
rect 174 601 176 603
rect 179 601 181 603
rect 184 601 186 603
rect 189 601 191 603
rect 194 601 196 603
rect 199 601 201 603
rect 204 601 206 603
rect 209 601 211 603
rect 214 601 216 603
rect 219 601 221 603
rect 224 601 226 603
rect 229 601 231 603
rect 234 601 236 603
rect 239 601 241 603
rect 244 601 246 603
rect 249 601 251 603
rect 254 601 256 603
rect 259 601 261 603
rect 264 601 266 603
rect 269 601 271 603
rect 274 601 276 603
rect 24 591 26 593
rect 29 591 31 593
rect 34 591 36 593
rect 39 591 41 593
rect 44 591 46 593
rect 49 591 51 593
rect 54 591 56 593
rect 59 591 61 593
rect 64 591 66 593
rect 69 591 71 593
rect 74 591 76 593
rect 79 591 81 593
rect 84 591 86 593
rect 89 591 91 593
rect 94 591 96 593
rect 99 591 101 593
rect 104 591 106 593
rect 109 591 111 593
rect 114 591 116 593
rect 119 591 121 593
rect 124 591 126 593
rect 129 591 131 593
rect 134 591 136 593
rect 139 591 141 593
rect 144 591 146 593
rect 149 591 151 593
rect 154 591 156 593
rect 159 591 161 593
rect 164 591 166 593
rect 169 591 171 593
rect 174 591 176 593
rect 179 591 181 593
rect 184 591 186 593
rect 189 591 191 593
rect 194 591 196 593
rect 199 591 201 593
rect 204 591 206 593
rect 209 591 211 593
rect 214 591 216 593
rect 219 591 221 593
rect 224 591 226 593
rect 229 591 231 593
rect 234 591 236 593
rect 239 591 241 593
rect 244 591 246 593
rect 249 591 251 593
rect 254 591 256 593
rect 259 591 261 593
rect 264 591 266 593
rect 269 591 271 593
rect 274 591 276 593
rect 24 581 26 583
rect 29 581 31 583
rect 34 581 36 583
rect 39 581 41 583
rect 44 581 46 583
rect 49 581 51 583
rect 54 581 56 583
rect 59 581 61 583
rect 64 581 66 583
rect 69 581 71 583
rect 74 581 76 583
rect 79 581 81 583
rect 84 581 86 583
rect 89 581 91 583
rect 94 581 96 583
rect 99 581 101 583
rect 104 581 106 583
rect 109 581 111 583
rect 114 581 116 583
rect 119 581 121 583
rect 124 581 126 583
rect 129 581 131 583
rect 134 581 136 583
rect 139 581 141 583
rect 144 581 146 583
rect 149 581 151 583
rect 154 581 156 583
rect 159 581 161 583
rect 164 581 166 583
rect 169 581 171 583
rect 174 581 176 583
rect 179 581 181 583
rect 184 581 186 583
rect 189 581 191 583
rect 194 581 196 583
rect 199 581 201 583
rect 204 581 206 583
rect 209 581 211 583
rect 214 581 216 583
rect 219 581 221 583
rect 224 581 226 583
rect 229 581 231 583
rect 234 581 236 583
rect 239 581 241 583
rect 244 581 246 583
rect 249 581 251 583
rect 254 581 256 583
rect 259 581 261 583
rect 264 581 266 583
rect 269 581 271 583
rect 274 581 276 583
rect 24 571 26 573
rect 29 571 31 573
rect 34 571 36 573
rect 39 571 41 573
rect 44 571 46 573
rect 49 571 51 573
rect 54 571 56 573
rect 59 571 61 573
rect 64 571 66 573
rect 69 571 71 573
rect 74 571 76 573
rect 79 571 81 573
rect 84 571 86 573
rect 89 571 91 573
rect 94 571 96 573
rect 99 571 101 573
rect 104 571 106 573
rect 109 571 111 573
rect 114 571 116 573
rect 119 571 121 573
rect 124 571 126 573
rect 129 571 131 573
rect 134 571 136 573
rect 139 571 141 573
rect 144 571 146 573
rect 149 571 151 573
rect 154 571 156 573
rect 159 571 161 573
rect 164 571 166 573
rect 169 571 171 573
rect 174 571 176 573
rect 179 571 181 573
rect 184 571 186 573
rect 189 571 191 573
rect 194 571 196 573
rect 199 571 201 573
rect 204 571 206 573
rect 209 571 211 573
rect 214 571 216 573
rect 219 571 221 573
rect 224 571 226 573
rect 229 571 231 573
rect 234 571 236 573
rect 239 571 241 573
rect 244 571 246 573
rect 249 571 251 573
rect 254 571 256 573
rect 259 571 261 573
rect 264 571 266 573
rect 269 571 271 573
rect 274 571 276 573
rect 24 561 26 563
rect 29 561 31 563
rect 34 561 36 563
rect 39 561 41 563
rect 44 561 46 563
rect 49 561 51 563
rect 54 561 56 563
rect 59 561 61 563
rect 64 561 66 563
rect 69 561 71 563
rect 74 561 76 563
rect 79 561 81 563
rect 84 561 86 563
rect 89 561 91 563
rect 94 561 96 563
rect 99 561 101 563
rect 104 561 106 563
rect 109 561 111 563
rect 114 561 116 563
rect 119 561 121 563
rect 124 561 126 563
rect 129 561 131 563
rect 134 561 136 563
rect 139 561 141 563
rect 144 561 146 563
rect 149 561 151 563
rect 154 561 156 563
rect 159 561 161 563
rect 164 561 166 563
rect 169 561 171 563
rect 174 561 176 563
rect 179 561 181 563
rect 184 561 186 563
rect 189 561 191 563
rect 194 561 196 563
rect 199 561 201 563
rect 204 561 206 563
rect 209 561 211 563
rect 214 561 216 563
rect 219 561 221 563
rect 224 561 226 563
rect 229 561 231 563
rect 234 561 236 563
rect 239 561 241 563
rect 244 561 246 563
rect 249 561 251 563
rect 254 561 256 563
rect 259 561 261 563
rect 264 561 266 563
rect 269 561 271 563
rect 274 561 276 563
rect 24 551 26 553
rect 29 551 31 553
rect 34 551 36 553
rect 39 551 41 553
rect 44 551 46 553
rect 49 551 51 553
rect 54 551 56 553
rect 59 551 61 553
rect 64 551 66 553
rect 69 551 71 553
rect 74 551 76 553
rect 79 551 81 553
rect 84 551 86 553
rect 89 551 91 553
rect 94 551 96 553
rect 99 551 101 553
rect 104 551 106 553
rect 109 551 111 553
rect 114 551 116 553
rect 119 551 121 553
rect 124 551 126 553
rect 129 551 131 553
rect 134 551 136 553
rect 139 551 141 553
rect 144 551 146 553
rect 149 551 151 553
rect 154 551 156 553
rect 159 551 161 553
rect 164 551 166 553
rect 169 551 171 553
rect 174 551 176 553
rect 179 551 181 553
rect 184 551 186 553
rect 189 551 191 553
rect 194 551 196 553
rect 199 551 201 553
rect 204 551 206 553
rect 209 551 211 553
rect 214 551 216 553
rect 219 551 221 553
rect 224 551 226 553
rect 229 551 231 553
rect 234 551 236 553
rect 239 551 241 553
rect 244 551 246 553
rect 249 551 251 553
rect 254 551 256 553
rect 259 551 261 553
rect 264 551 266 553
rect 269 551 271 553
rect 274 551 276 553
rect 24 541 26 543
rect 29 541 31 543
rect 34 541 36 543
rect 39 541 41 543
rect 44 541 46 543
rect 49 541 51 543
rect 54 541 56 543
rect 59 541 61 543
rect 64 541 66 543
rect 69 541 71 543
rect 74 541 76 543
rect 79 541 81 543
rect 84 541 86 543
rect 89 541 91 543
rect 94 541 96 543
rect 99 541 101 543
rect 104 541 106 543
rect 109 541 111 543
rect 114 541 116 543
rect 119 541 121 543
rect 124 541 126 543
rect 129 541 131 543
rect 134 541 136 543
rect 139 541 141 543
rect 144 541 146 543
rect 149 541 151 543
rect 154 541 156 543
rect 159 541 161 543
rect 164 541 166 543
rect 169 541 171 543
rect 174 541 176 543
rect 179 541 181 543
rect 184 541 186 543
rect 189 541 191 543
rect 194 541 196 543
rect 199 541 201 543
rect 204 541 206 543
rect 209 541 211 543
rect 214 541 216 543
rect 219 541 221 543
rect 224 541 226 543
rect 229 541 231 543
rect 234 541 236 543
rect 239 541 241 543
rect 244 541 246 543
rect 249 541 251 543
rect 254 541 256 543
rect 259 541 261 543
rect 264 541 266 543
rect 269 541 271 543
rect 274 541 276 543
rect 24 531 26 533
rect 29 531 31 533
rect 34 531 36 533
rect 39 531 41 533
rect 44 531 46 533
rect 49 531 51 533
rect 54 531 56 533
rect 59 531 61 533
rect 64 531 66 533
rect 69 531 71 533
rect 74 531 76 533
rect 79 531 81 533
rect 84 531 86 533
rect 89 531 91 533
rect 94 531 96 533
rect 99 531 101 533
rect 104 531 106 533
rect 109 531 111 533
rect 114 531 116 533
rect 119 531 121 533
rect 124 531 126 533
rect 129 531 131 533
rect 134 531 136 533
rect 139 531 141 533
rect 144 531 146 533
rect 149 531 151 533
rect 154 531 156 533
rect 159 531 161 533
rect 164 531 166 533
rect 169 531 171 533
rect 174 531 176 533
rect 179 531 181 533
rect 184 531 186 533
rect 189 531 191 533
rect 194 531 196 533
rect 199 531 201 533
rect 204 531 206 533
rect 209 531 211 533
rect 214 531 216 533
rect 219 531 221 533
rect 224 531 226 533
rect 229 531 231 533
rect 234 531 236 533
rect 239 531 241 533
rect 244 531 246 533
rect 249 531 251 533
rect 254 531 256 533
rect 259 531 261 533
rect 264 531 266 533
rect 269 531 271 533
rect 274 531 276 533
rect 24 521 26 523
rect 29 521 31 523
rect 34 521 36 523
rect 39 521 41 523
rect 44 521 46 523
rect 49 521 51 523
rect 54 521 56 523
rect 59 521 61 523
rect 64 521 66 523
rect 69 521 71 523
rect 74 521 76 523
rect 79 521 81 523
rect 84 521 86 523
rect 89 521 91 523
rect 94 521 96 523
rect 99 521 101 523
rect 104 521 106 523
rect 109 521 111 523
rect 114 521 116 523
rect 119 521 121 523
rect 124 521 126 523
rect 129 521 131 523
rect 134 521 136 523
rect 139 521 141 523
rect 144 521 146 523
rect 149 521 151 523
rect 154 521 156 523
rect 159 521 161 523
rect 164 521 166 523
rect 169 521 171 523
rect 174 521 176 523
rect 179 521 181 523
rect 184 521 186 523
rect 189 521 191 523
rect 194 521 196 523
rect 199 521 201 523
rect 204 521 206 523
rect 209 521 211 523
rect 214 521 216 523
rect 219 521 221 523
rect 224 521 226 523
rect 229 521 231 523
rect 234 521 236 523
rect 239 521 241 523
rect 244 521 246 523
rect 249 521 251 523
rect 254 521 256 523
rect 259 521 261 523
rect 264 521 266 523
rect 269 521 271 523
rect 274 521 276 523
rect 24 511 26 513
rect 29 511 31 513
rect 34 511 36 513
rect 39 511 41 513
rect 44 511 46 513
rect 49 511 51 513
rect 54 511 56 513
rect 59 511 61 513
rect 64 511 66 513
rect 69 511 71 513
rect 74 511 76 513
rect 79 511 81 513
rect 84 511 86 513
rect 89 511 91 513
rect 94 511 96 513
rect 99 511 101 513
rect 104 511 106 513
rect 109 511 111 513
rect 114 511 116 513
rect 119 511 121 513
rect 124 511 126 513
rect 129 511 131 513
rect 134 511 136 513
rect 139 511 141 513
rect 144 511 146 513
rect 149 511 151 513
rect 154 511 156 513
rect 159 511 161 513
rect 164 511 166 513
rect 169 511 171 513
rect 174 511 176 513
rect 179 511 181 513
rect 184 511 186 513
rect 189 511 191 513
rect 194 511 196 513
rect 199 511 201 513
rect 204 511 206 513
rect 209 511 211 513
rect 214 511 216 513
rect 219 511 221 513
rect 224 511 226 513
rect 229 511 231 513
rect 234 511 236 513
rect 239 511 241 513
rect 244 511 246 513
rect 249 511 251 513
rect 254 511 256 513
rect 259 511 261 513
rect 264 511 266 513
rect 269 511 271 513
rect 274 511 276 513
rect 24 501 26 503
rect 29 501 31 503
rect 34 501 36 503
rect 39 501 41 503
rect 44 501 46 503
rect 49 501 51 503
rect 54 501 56 503
rect 59 501 61 503
rect 64 501 66 503
rect 69 501 71 503
rect 74 501 76 503
rect 79 501 81 503
rect 84 501 86 503
rect 89 501 91 503
rect 94 501 96 503
rect 99 501 101 503
rect 104 501 106 503
rect 109 501 111 503
rect 114 501 116 503
rect 119 501 121 503
rect 124 501 126 503
rect 129 501 131 503
rect 134 501 136 503
rect 139 501 141 503
rect 144 501 146 503
rect 149 501 151 503
rect 154 501 156 503
rect 159 501 161 503
rect 164 501 166 503
rect 169 501 171 503
rect 174 501 176 503
rect 179 501 181 503
rect 184 501 186 503
rect 189 501 191 503
rect 194 501 196 503
rect 199 501 201 503
rect 204 501 206 503
rect 209 501 211 503
rect 214 501 216 503
rect 219 501 221 503
rect 224 501 226 503
rect 229 501 231 503
rect 234 501 236 503
rect 239 501 241 503
rect 244 501 246 503
rect 249 501 251 503
rect 254 501 256 503
rect 259 501 261 503
rect 264 501 266 503
rect 269 501 271 503
rect 274 501 276 503
rect 24 491 26 493
rect 29 491 31 493
rect 34 491 36 493
rect 39 491 41 493
rect 44 491 46 493
rect 49 491 51 493
rect 54 491 56 493
rect 59 491 61 493
rect 64 491 66 493
rect 69 491 71 493
rect 74 491 76 493
rect 79 491 81 493
rect 84 491 86 493
rect 89 491 91 493
rect 94 491 96 493
rect 99 491 101 493
rect 104 491 106 493
rect 109 491 111 493
rect 114 491 116 493
rect 119 491 121 493
rect 124 491 126 493
rect 129 491 131 493
rect 134 491 136 493
rect 139 491 141 493
rect 144 491 146 493
rect 149 491 151 493
rect 154 491 156 493
rect 159 491 161 493
rect 164 491 166 493
rect 169 491 171 493
rect 174 491 176 493
rect 179 491 181 493
rect 184 491 186 493
rect 189 491 191 493
rect 194 491 196 493
rect 199 491 201 493
rect 204 491 206 493
rect 209 491 211 493
rect 214 491 216 493
rect 219 491 221 493
rect 224 491 226 493
rect 229 491 231 493
rect 234 491 236 493
rect 239 491 241 493
rect 244 491 246 493
rect 249 491 251 493
rect 254 491 256 493
rect 259 491 261 493
rect 264 491 266 493
rect 269 491 271 493
rect 274 491 276 493
rect 24 481 26 483
rect 29 481 31 483
rect 34 481 36 483
rect 39 481 41 483
rect 44 481 46 483
rect 49 481 51 483
rect 54 481 56 483
rect 59 481 61 483
rect 64 481 66 483
rect 69 481 71 483
rect 74 481 76 483
rect 79 481 81 483
rect 84 481 86 483
rect 89 481 91 483
rect 94 481 96 483
rect 99 481 101 483
rect 104 481 106 483
rect 109 481 111 483
rect 114 481 116 483
rect 119 481 121 483
rect 124 481 126 483
rect 129 481 131 483
rect 134 481 136 483
rect 139 481 141 483
rect 144 481 146 483
rect 149 481 151 483
rect 154 481 156 483
rect 159 481 161 483
rect 164 481 166 483
rect 169 481 171 483
rect 174 481 176 483
rect 179 481 181 483
rect 184 481 186 483
rect 189 481 191 483
rect 194 481 196 483
rect 199 481 201 483
rect 204 481 206 483
rect 209 481 211 483
rect 214 481 216 483
rect 219 481 221 483
rect 224 481 226 483
rect 229 481 231 483
rect 234 481 236 483
rect 239 481 241 483
rect 244 481 246 483
rect 249 481 251 483
rect 254 481 256 483
rect 259 481 261 483
rect 264 481 266 483
rect 269 481 271 483
rect 274 481 276 483
rect 24 471 26 473
rect 29 471 31 473
rect 34 471 36 473
rect 39 471 41 473
rect 44 471 46 473
rect 49 471 51 473
rect 54 471 56 473
rect 59 471 61 473
rect 64 471 66 473
rect 69 471 71 473
rect 74 471 76 473
rect 79 471 81 473
rect 84 471 86 473
rect 89 471 91 473
rect 94 471 96 473
rect 99 471 101 473
rect 104 471 106 473
rect 109 471 111 473
rect 114 471 116 473
rect 119 471 121 473
rect 124 471 126 473
rect 129 471 131 473
rect 134 471 136 473
rect 139 471 141 473
rect 144 471 146 473
rect 149 471 151 473
rect 154 471 156 473
rect 159 471 161 473
rect 164 471 166 473
rect 169 471 171 473
rect 174 471 176 473
rect 179 471 181 473
rect 184 471 186 473
rect 189 471 191 473
rect 194 471 196 473
rect 199 471 201 473
rect 204 471 206 473
rect 209 471 211 473
rect 214 471 216 473
rect 219 471 221 473
rect 224 471 226 473
rect 229 471 231 473
rect 234 471 236 473
rect 239 471 241 473
rect 244 471 246 473
rect 249 471 251 473
rect 254 471 256 473
rect 259 471 261 473
rect 264 471 266 473
rect 269 471 271 473
rect 274 471 276 473
rect 24 461 26 463
rect 29 461 31 463
rect 34 461 36 463
rect 39 461 41 463
rect 44 461 46 463
rect 49 461 51 463
rect 54 461 56 463
rect 59 461 61 463
rect 64 461 66 463
rect 69 461 71 463
rect 74 461 76 463
rect 79 461 81 463
rect 84 461 86 463
rect 89 461 91 463
rect 94 461 96 463
rect 99 461 101 463
rect 104 461 106 463
rect 109 461 111 463
rect 114 461 116 463
rect 119 461 121 463
rect 124 461 126 463
rect 129 461 131 463
rect 134 461 136 463
rect 139 461 141 463
rect 144 461 146 463
rect 149 461 151 463
rect 154 461 156 463
rect 159 461 161 463
rect 164 461 166 463
rect 169 461 171 463
rect 174 461 176 463
rect 179 461 181 463
rect 184 461 186 463
rect 189 461 191 463
rect 194 461 196 463
rect 199 461 201 463
rect 204 461 206 463
rect 209 461 211 463
rect 214 461 216 463
rect 219 461 221 463
rect 224 461 226 463
rect 229 461 231 463
rect 234 461 236 463
rect 239 461 241 463
rect 244 461 246 463
rect 249 461 251 463
rect 254 461 256 463
rect 259 461 261 463
rect 264 461 266 463
rect 269 461 271 463
rect 274 461 276 463
rect 24 451 26 453
rect 29 451 31 453
rect 34 451 36 453
rect 39 451 41 453
rect 44 451 46 453
rect 49 451 51 453
rect 54 451 56 453
rect 59 451 61 453
rect 64 451 66 453
rect 69 451 71 453
rect 74 451 76 453
rect 79 451 81 453
rect 84 451 86 453
rect 89 451 91 453
rect 94 451 96 453
rect 99 451 101 453
rect 104 451 106 453
rect 109 451 111 453
rect 114 451 116 453
rect 119 451 121 453
rect 124 451 126 453
rect 129 451 131 453
rect 134 451 136 453
rect 139 451 141 453
rect 144 451 146 453
rect 149 451 151 453
rect 154 451 156 453
rect 159 451 161 453
rect 164 451 166 453
rect 169 451 171 453
rect 174 451 176 453
rect 179 451 181 453
rect 184 451 186 453
rect 189 451 191 453
rect 194 451 196 453
rect 199 451 201 453
rect 204 451 206 453
rect 209 451 211 453
rect 214 451 216 453
rect 219 451 221 453
rect 224 451 226 453
rect 229 451 231 453
rect 234 451 236 453
rect 239 451 241 453
rect 244 451 246 453
rect 249 451 251 453
rect 254 451 256 453
rect 259 451 261 453
rect 264 451 266 453
rect 269 451 271 453
rect 274 451 276 453
rect 24 441 26 443
rect 29 441 31 443
rect 34 441 36 443
rect 39 441 41 443
rect 44 441 46 443
rect 49 441 51 443
rect 54 441 56 443
rect 59 441 61 443
rect 64 441 66 443
rect 69 441 71 443
rect 74 441 76 443
rect 79 441 81 443
rect 84 441 86 443
rect 89 441 91 443
rect 94 441 96 443
rect 99 441 101 443
rect 104 441 106 443
rect 109 441 111 443
rect 114 441 116 443
rect 119 441 121 443
rect 124 441 126 443
rect 129 441 131 443
rect 134 441 136 443
rect 139 441 141 443
rect 144 441 146 443
rect 149 441 151 443
rect 154 441 156 443
rect 159 441 161 443
rect 164 441 166 443
rect 169 441 171 443
rect 174 441 176 443
rect 179 441 181 443
rect 184 441 186 443
rect 189 441 191 443
rect 194 441 196 443
rect 199 441 201 443
rect 204 441 206 443
rect 209 441 211 443
rect 214 441 216 443
rect 219 441 221 443
rect 224 441 226 443
rect 229 441 231 443
rect 234 441 236 443
rect 239 441 241 443
rect 244 441 246 443
rect 249 441 251 443
rect 254 441 256 443
rect 259 441 261 443
rect 264 441 266 443
rect 269 441 271 443
rect 274 441 276 443
rect 3 415 5 417
rect 8 415 10 417
rect 13 415 15 417
rect 18 415 20 417
rect 23 415 25 417
rect 28 415 30 417
rect 33 415 35 417
rect 38 415 40 417
rect 43 415 45 417
rect 48 415 50 417
rect 53 415 55 417
rect 58 415 60 417
rect 63 415 65 417
rect 68 415 70 417
rect 73 415 75 417
rect 78 415 80 417
rect 83 415 85 417
rect 88 415 90 417
rect 93 415 95 417
rect 144 410 146 412
rect 149 410 151 412
rect 154 410 156 412
rect 205 410 207 412
rect 210 410 212 412
rect 215 410 217 412
rect 220 410 222 412
rect 225 410 227 412
rect 230 410 232 412
rect 235 410 237 412
rect 240 410 242 412
rect 245 410 247 412
rect 250 410 252 412
rect 255 410 257 412
rect 260 410 262 412
rect 265 410 267 412
rect 270 410 272 412
rect 275 410 277 412
rect 280 410 282 412
rect 285 410 287 412
rect 290 410 292 412
rect 295 410 297 412
rect 3 405 5 407
rect 8 405 10 407
rect 13 405 15 407
rect 18 405 20 407
rect 23 405 25 407
rect 28 405 30 407
rect 33 405 35 407
rect 38 405 40 407
rect 43 405 45 407
rect 48 405 50 407
rect 53 405 55 407
rect 58 405 60 407
rect 63 405 65 407
rect 68 405 70 407
rect 73 405 75 407
rect 78 405 80 407
rect 83 405 85 407
rect 88 405 90 407
rect 93 405 95 407
rect 144 400 146 402
rect 149 400 151 402
rect 154 400 156 402
rect 205 400 207 402
rect 210 400 212 402
rect 215 400 217 402
rect 220 400 222 402
rect 225 400 227 402
rect 230 400 232 402
rect 235 400 237 402
rect 240 400 242 402
rect 245 400 247 402
rect 250 400 252 402
rect 255 400 257 402
rect 260 400 262 402
rect 265 400 267 402
rect 270 400 272 402
rect 275 400 277 402
rect 280 400 282 402
rect 285 400 287 402
rect 290 400 292 402
rect 295 400 297 402
rect 3 395 5 397
rect 8 395 10 397
rect 13 395 15 397
rect 18 395 20 397
rect 23 395 25 397
rect 28 395 30 397
rect 33 395 35 397
rect 38 395 40 397
rect 43 395 45 397
rect 48 395 50 397
rect 53 395 55 397
rect 58 395 60 397
rect 63 395 65 397
rect 68 395 70 397
rect 73 395 75 397
rect 78 395 80 397
rect 83 395 85 397
rect 88 395 90 397
rect 93 395 95 397
rect 144 390 146 392
rect 149 390 151 392
rect 154 390 156 392
rect 205 390 207 392
rect 210 390 212 392
rect 215 390 217 392
rect 220 390 222 392
rect 225 390 227 392
rect 230 390 232 392
rect 235 390 237 392
rect 240 390 242 392
rect 245 390 247 392
rect 250 390 252 392
rect 255 390 257 392
rect 260 390 262 392
rect 265 390 267 392
rect 270 390 272 392
rect 275 390 277 392
rect 280 390 282 392
rect 285 390 287 392
rect 290 390 292 392
rect 295 390 297 392
rect 3 385 5 387
rect 8 385 10 387
rect 13 385 15 387
rect 18 385 20 387
rect 23 385 25 387
rect 28 385 30 387
rect 33 385 35 387
rect 38 385 40 387
rect 43 385 45 387
rect 48 385 50 387
rect 53 385 55 387
rect 58 385 60 387
rect 63 385 65 387
rect 68 385 70 387
rect 73 385 75 387
rect 78 385 80 387
rect 83 385 85 387
rect 88 385 90 387
rect 93 385 95 387
rect 144 380 146 382
rect 149 380 151 382
rect 154 380 156 382
rect 205 380 207 382
rect 210 380 212 382
rect 215 380 217 382
rect 220 380 222 382
rect 225 380 227 382
rect 230 380 232 382
rect 235 380 237 382
rect 240 380 242 382
rect 245 380 247 382
rect 250 380 252 382
rect 255 380 257 382
rect 260 380 262 382
rect 265 380 267 382
rect 270 380 272 382
rect 275 380 277 382
rect 280 380 282 382
rect 285 380 287 382
rect 290 380 292 382
rect 295 380 297 382
rect 3 375 5 377
rect 8 375 10 377
rect 13 375 15 377
rect 18 375 20 377
rect 23 375 25 377
rect 28 375 30 377
rect 33 375 35 377
rect 38 375 40 377
rect 43 375 45 377
rect 48 375 50 377
rect 53 375 55 377
rect 58 375 60 377
rect 63 375 65 377
rect 68 375 70 377
rect 73 375 75 377
rect 78 375 80 377
rect 83 375 85 377
rect 88 375 90 377
rect 93 375 95 377
rect 144 370 146 372
rect 149 370 151 372
rect 154 370 156 372
rect 205 370 207 372
rect 210 370 212 372
rect 215 370 217 372
rect 220 370 222 372
rect 225 370 227 372
rect 230 370 232 372
rect 235 370 237 372
rect 240 370 242 372
rect 245 370 247 372
rect 250 370 252 372
rect 255 370 257 372
rect 260 370 262 372
rect 265 370 267 372
rect 270 370 272 372
rect 275 370 277 372
rect 280 370 282 372
rect 285 370 287 372
rect 290 370 292 372
rect 295 370 297 372
rect 3 365 5 367
rect 8 365 10 367
rect 13 365 15 367
rect 18 365 20 367
rect 23 365 25 367
rect 28 365 30 367
rect 33 365 35 367
rect 38 365 40 367
rect 43 365 45 367
rect 48 365 50 367
rect 53 365 55 367
rect 58 365 60 367
rect 63 365 65 367
rect 68 365 70 367
rect 73 365 75 367
rect 78 365 80 367
rect 83 365 85 367
rect 88 365 90 367
rect 93 365 95 367
rect 144 360 146 362
rect 149 360 151 362
rect 154 360 156 362
rect 205 360 207 362
rect 210 360 212 362
rect 215 360 217 362
rect 220 360 222 362
rect 225 360 227 362
rect 230 360 232 362
rect 235 360 237 362
rect 240 360 242 362
rect 245 360 247 362
rect 250 360 252 362
rect 255 360 257 362
rect 260 360 262 362
rect 265 360 267 362
rect 270 360 272 362
rect 275 360 277 362
rect 280 360 282 362
rect 285 360 287 362
rect 290 360 292 362
rect 295 360 297 362
rect 3 355 5 357
rect 8 355 10 357
rect 13 355 15 357
rect 18 355 20 357
rect 23 355 25 357
rect 28 355 30 357
rect 33 355 35 357
rect 38 355 40 357
rect 43 355 45 357
rect 48 355 50 357
rect 53 355 55 357
rect 58 355 60 357
rect 63 355 65 357
rect 68 355 70 357
rect 73 355 75 357
rect 78 355 80 357
rect 83 355 85 357
rect 88 355 90 357
rect 93 355 95 357
rect 3 350 5 352
rect 8 350 10 352
rect 13 350 15 352
rect 18 350 20 352
rect 23 350 25 352
rect 28 350 30 352
rect 33 350 35 352
rect 38 350 40 352
rect 43 350 45 352
rect 48 350 50 352
rect 53 350 55 352
rect 58 350 60 352
rect 63 350 65 352
rect 68 350 70 352
rect 73 350 75 352
rect 78 350 80 352
rect 83 350 85 352
rect 88 350 90 352
rect 93 350 95 352
rect 144 350 146 352
rect 149 350 151 352
rect 154 350 156 352
rect 205 350 207 352
rect 210 350 212 352
rect 215 350 217 352
rect 220 350 222 352
rect 225 350 227 352
rect 230 350 232 352
rect 235 350 237 352
rect 240 350 242 352
rect 245 350 247 352
rect 250 350 252 352
rect 255 350 257 352
rect 260 350 262 352
rect 265 350 267 352
rect 270 350 272 352
rect 275 350 277 352
rect 280 350 282 352
rect 285 350 287 352
rect 290 350 292 352
rect 295 350 297 352
rect 4 318 6 320
rect 9 318 11 320
rect 14 318 16 320
rect 19 318 21 320
rect 24 318 26 320
rect 29 318 31 320
rect 34 318 36 320
rect 39 318 41 320
rect 44 318 46 320
rect 49 318 51 320
rect 54 318 56 320
rect 59 318 61 320
rect 64 318 66 320
rect 69 318 71 320
rect 74 318 76 320
rect 79 318 81 320
rect 84 318 86 320
rect 89 318 91 320
rect 94 318 96 320
rect 99 318 101 320
rect 104 318 106 320
rect 109 318 111 320
rect 114 318 116 320
rect 119 318 121 320
rect 124 318 126 320
rect 129 318 131 320
rect 134 318 136 320
rect 139 318 141 320
rect 144 318 146 320
rect 149 318 151 320
rect 154 318 156 320
rect 159 318 161 320
rect 164 318 166 320
rect 169 318 171 320
rect 174 318 176 320
rect 179 318 181 320
rect 184 318 186 320
rect 189 318 191 320
rect 194 318 196 320
rect 199 318 201 320
rect 204 318 206 320
rect 209 318 211 320
rect 214 318 216 320
rect 219 318 221 320
rect 224 318 226 320
rect 229 318 231 320
rect 234 318 236 320
rect 239 318 241 320
rect 244 318 246 320
rect 249 318 251 320
rect 254 318 256 320
rect 259 318 261 320
rect 264 318 266 320
rect 269 318 271 320
rect 274 318 276 320
rect 279 318 281 320
rect 284 318 286 320
rect 289 318 291 320
rect 294 318 296 320
rect 4 308 6 310
rect 9 308 11 310
rect 14 308 16 310
rect 19 308 21 310
rect 24 308 26 310
rect 29 308 31 310
rect 34 308 36 310
rect 39 308 41 310
rect 44 308 46 310
rect 49 308 51 310
rect 54 308 56 310
rect 59 308 61 310
rect 64 308 66 310
rect 69 308 71 310
rect 74 308 76 310
rect 79 308 81 310
rect 84 308 86 310
rect 89 308 91 310
rect 94 308 96 310
rect 99 308 101 310
rect 104 308 106 310
rect 109 308 111 310
rect 114 308 116 310
rect 119 308 121 310
rect 124 308 126 310
rect 129 308 131 310
rect 134 308 136 310
rect 139 308 141 310
rect 144 308 146 310
rect 149 308 151 310
rect 154 308 156 310
rect 159 308 161 310
rect 164 308 166 310
rect 169 308 171 310
rect 174 308 176 310
rect 179 308 181 310
rect 184 308 186 310
rect 189 308 191 310
rect 194 308 196 310
rect 199 308 201 310
rect 204 308 206 310
rect 209 308 211 310
rect 214 308 216 310
rect 219 308 221 310
rect 224 308 226 310
rect 229 308 231 310
rect 234 308 236 310
rect 239 308 241 310
rect 244 308 246 310
rect 249 308 251 310
rect 254 308 256 310
rect 259 308 261 310
rect 264 308 266 310
rect 269 308 271 310
rect 274 308 276 310
rect 279 308 281 310
rect 284 308 286 310
rect 289 308 291 310
rect 294 308 296 310
rect 4 298 6 300
rect 9 298 11 300
rect 14 298 16 300
rect 19 298 21 300
rect 24 298 26 300
rect 29 298 31 300
rect 34 298 36 300
rect 39 298 41 300
rect 44 298 46 300
rect 49 298 51 300
rect 54 298 56 300
rect 59 298 61 300
rect 64 298 66 300
rect 69 298 71 300
rect 74 298 76 300
rect 79 298 81 300
rect 84 298 86 300
rect 89 298 91 300
rect 94 298 96 300
rect 99 298 101 300
rect 104 298 106 300
rect 109 298 111 300
rect 114 298 116 300
rect 119 298 121 300
rect 124 298 126 300
rect 129 298 131 300
rect 134 298 136 300
rect 139 298 141 300
rect 144 298 146 300
rect 149 298 151 300
rect 154 298 156 300
rect 159 298 161 300
rect 164 298 166 300
rect 169 298 171 300
rect 174 298 176 300
rect 179 298 181 300
rect 184 298 186 300
rect 189 298 191 300
rect 194 298 196 300
rect 199 298 201 300
rect 204 298 206 300
rect 209 298 211 300
rect 214 298 216 300
rect 219 298 221 300
rect 224 298 226 300
rect 229 298 231 300
rect 234 298 236 300
rect 239 298 241 300
rect 244 298 246 300
rect 249 298 251 300
rect 254 298 256 300
rect 259 298 261 300
rect 264 298 266 300
rect 269 298 271 300
rect 274 298 276 300
rect 279 298 281 300
rect 284 298 286 300
rect 289 298 291 300
rect 294 298 296 300
rect 4 288 6 290
rect 9 288 11 290
rect 14 288 16 290
rect 19 288 21 290
rect 24 288 26 290
rect 29 288 31 290
rect 34 288 36 290
rect 39 288 41 290
rect 44 288 46 290
rect 49 288 51 290
rect 54 288 56 290
rect 59 288 61 290
rect 64 288 66 290
rect 69 288 71 290
rect 74 288 76 290
rect 79 288 81 290
rect 84 288 86 290
rect 89 288 91 290
rect 94 288 96 290
rect 99 288 101 290
rect 104 288 106 290
rect 109 288 111 290
rect 114 288 116 290
rect 119 288 121 290
rect 124 288 126 290
rect 129 288 131 290
rect 134 288 136 290
rect 139 288 141 290
rect 144 288 146 290
rect 149 288 151 290
rect 154 288 156 290
rect 159 288 161 290
rect 164 288 166 290
rect 169 288 171 290
rect 174 288 176 290
rect 179 288 181 290
rect 184 288 186 290
rect 189 288 191 290
rect 194 288 196 290
rect 199 288 201 290
rect 204 288 206 290
rect 209 288 211 290
rect 214 288 216 290
rect 219 288 221 290
rect 224 288 226 290
rect 229 288 231 290
rect 234 288 236 290
rect 239 288 241 290
rect 244 288 246 290
rect 249 288 251 290
rect 254 288 256 290
rect 259 288 261 290
rect 264 288 266 290
rect 269 288 271 290
rect 274 288 276 290
rect 279 288 281 290
rect 284 288 286 290
rect 289 288 291 290
rect 294 288 296 290
rect 4 278 6 280
rect 9 278 11 280
rect 14 278 16 280
rect 19 278 21 280
rect 24 278 26 280
rect 29 278 31 280
rect 34 278 36 280
rect 39 278 41 280
rect 44 278 46 280
rect 49 278 51 280
rect 54 278 56 280
rect 59 278 61 280
rect 64 278 66 280
rect 69 278 71 280
rect 74 278 76 280
rect 79 278 81 280
rect 84 278 86 280
rect 89 278 91 280
rect 94 278 96 280
rect 99 278 101 280
rect 104 278 106 280
rect 109 278 111 280
rect 114 278 116 280
rect 119 278 121 280
rect 124 278 126 280
rect 129 278 131 280
rect 134 278 136 280
rect 139 278 141 280
rect 144 278 146 280
rect 149 278 151 280
rect 154 278 156 280
rect 159 278 161 280
rect 164 278 166 280
rect 169 278 171 280
rect 174 278 176 280
rect 179 278 181 280
rect 184 278 186 280
rect 189 278 191 280
rect 194 278 196 280
rect 199 278 201 280
rect 204 278 206 280
rect 209 278 211 280
rect 214 278 216 280
rect 219 278 221 280
rect 224 278 226 280
rect 229 278 231 280
rect 234 278 236 280
rect 239 278 241 280
rect 244 278 246 280
rect 249 278 251 280
rect 254 278 256 280
rect 259 278 261 280
rect 264 278 266 280
rect 269 278 271 280
rect 274 278 276 280
rect 279 278 281 280
rect 284 278 286 280
rect 289 278 291 280
rect 294 278 296 280
rect 4 268 6 270
rect 9 268 11 270
rect 14 268 16 270
rect 19 268 21 270
rect 24 268 26 270
rect 29 268 31 270
rect 34 268 36 270
rect 39 268 41 270
rect 44 268 46 270
rect 49 268 51 270
rect 54 268 56 270
rect 59 268 61 270
rect 64 268 66 270
rect 69 268 71 270
rect 74 268 76 270
rect 79 268 81 270
rect 84 268 86 270
rect 89 268 91 270
rect 94 268 96 270
rect 99 268 101 270
rect 104 268 106 270
rect 109 268 111 270
rect 114 268 116 270
rect 119 268 121 270
rect 124 268 126 270
rect 129 268 131 270
rect 134 268 136 270
rect 139 268 141 270
rect 144 268 146 270
rect 149 268 151 270
rect 154 268 156 270
rect 159 268 161 270
rect 164 268 166 270
rect 169 268 171 270
rect 174 268 176 270
rect 179 268 181 270
rect 184 268 186 270
rect 189 268 191 270
rect 194 268 196 270
rect 199 268 201 270
rect 204 268 206 270
rect 209 268 211 270
rect 214 268 216 270
rect 219 268 221 270
rect 224 268 226 270
rect 229 268 231 270
rect 234 268 236 270
rect 239 268 241 270
rect 244 268 246 270
rect 249 268 251 270
rect 254 268 256 270
rect 259 268 261 270
rect 264 268 266 270
rect 269 268 271 270
rect 274 268 276 270
rect 279 268 281 270
rect 284 268 286 270
rect 289 268 291 270
rect 294 268 296 270
rect 9 258 11 260
rect 14 258 16 260
rect 19 258 21 260
rect 24 258 26 260
rect 29 258 31 260
rect 34 258 36 260
rect 39 258 41 260
rect 44 258 46 260
rect 49 258 51 260
rect 54 258 56 260
rect 59 258 61 260
rect 64 258 66 260
rect 69 258 71 260
rect 74 258 76 260
rect 79 258 81 260
rect 84 258 86 260
rect 89 258 91 260
rect 94 258 96 260
rect 99 258 101 260
rect 104 258 106 260
rect 109 258 111 260
rect 114 258 116 260
rect 119 258 121 260
rect 124 258 126 260
rect 129 258 131 260
rect 134 258 136 260
rect 139 258 141 260
rect 144 258 146 260
rect 149 258 151 260
rect 154 258 156 260
rect 159 258 161 260
rect 164 258 166 260
rect 169 258 171 260
rect 174 258 176 260
rect 179 258 181 260
rect 184 258 186 260
rect 189 258 191 260
rect 194 258 196 260
rect 199 258 201 260
rect 204 258 206 260
rect 209 258 211 260
rect 214 258 216 260
rect 219 258 221 260
rect 224 258 226 260
rect 229 258 231 260
rect 234 258 236 260
rect 239 258 241 260
rect 244 258 246 260
rect 249 258 251 260
rect 254 258 256 260
rect 259 258 261 260
rect 264 258 266 260
rect 269 258 271 260
rect 274 258 276 260
rect 279 258 281 260
rect 284 258 286 260
rect 289 258 291 260
rect 20 224 22 226
rect 146 223 148 225
rect 151 223 153 225
rect 273 224 275 226
rect 20 219 22 221
rect 273 219 275 221
rect 20 214 22 216
rect 146 215 148 217
rect 151 215 153 217
rect 273 214 275 216
rect 40 211 42 213
rect 45 211 47 213
rect 50 211 52 213
rect 58 211 60 213
rect 63 211 65 213
rect 68 211 70 213
rect 73 211 75 213
rect 78 211 80 213
rect 83 211 85 213
rect 88 211 90 213
rect 93 211 95 213
rect 205 211 207 213
rect 210 211 212 213
rect 215 211 217 213
rect 220 211 222 213
rect 225 211 227 213
rect 230 211 232 213
rect 235 211 237 213
rect 240 211 242 213
rect 248 211 250 213
rect 253 211 255 213
rect 258 211 260 213
rect 20 209 22 211
rect 273 209 275 211
rect 40 206 42 208
rect 45 206 47 208
rect 50 206 52 208
rect 146 207 148 209
rect 151 207 153 209
rect 248 206 250 208
rect 253 206 255 208
rect 258 206 260 208
rect 20 204 22 206
rect 273 204 275 206
rect 40 201 42 203
rect 45 201 47 203
rect 50 201 52 203
rect 248 201 250 203
rect 253 201 255 203
rect 258 201 260 203
rect 20 199 22 201
rect 273 199 275 201
rect 40 196 42 198
rect 45 196 47 198
rect 50 196 52 198
rect 248 196 250 198
rect 253 196 255 198
rect 258 196 260 198
rect 20 194 22 196
rect 273 194 275 196
rect 20 189 22 191
rect 40 190 42 192
rect 45 190 47 192
rect 50 190 52 192
rect 248 190 250 192
rect 253 190 255 192
rect 258 190 260 192
rect 273 189 275 191
rect 20 184 22 186
rect 40 185 42 187
rect 45 185 47 187
rect 50 185 52 187
rect 248 185 250 187
rect 253 185 255 187
rect 258 185 260 187
rect 273 184 275 186
rect 20 179 22 181
rect 40 180 42 182
rect 45 180 47 182
rect 50 180 52 182
rect 248 180 250 182
rect 253 180 255 182
rect 258 180 260 182
rect 273 179 275 181
rect 20 174 22 176
rect 40 175 42 177
rect 45 175 47 177
rect 50 175 52 177
rect 58 175 60 177
rect 63 175 65 177
rect 68 175 70 177
rect 73 175 75 177
rect 78 175 80 177
rect 83 175 85 177
rect 88 175 90 177
rect 93 175 95 177
rect 98 175 100 177
rect 103 175 105 177
rect 108 175 110 177
rect 113 175 115 177
rect 185 175 187 177
rect 190 175 192 177
rect 195 175 197 177
rect 200 175 202 177
rect 205 175 207 177
rect 210 175 212 177
rect 215 175 217 177
rect 220 175 222 177
rect 225 175 227 177
rect 230 175 232 177
rect 235 175 237 177
rect 240 175 242 177
rect 248 175 250 177
rect 253 175 255 177
rect 258 175 260 177
rect 273 174 275 176
rect 20 169 22 171
rect 273 169 275 171
rect 20 164 22 166
rect 273 164 275 166
rect 20 159 22 161
rect 273 159 275 161
rect 20 154 22 156
rect 273 154 275 156
rect 20 149 22 151
rect 273 149 275 151
rect 20 144 22 146
rect 40 145 42 147
rect 45 145 47 147
rect 50 145 52 147
rect 58 145 60 147
rect 63 145 65 147
rect 68 145 70 147
rect 73 145 75 147
rect 78 145 80 147
rect 83 145 85 147
rect 88 145 90 147
rect 93 145 95 147
rect 98 145 100 147
rect 103 145 105 147
rect 108 145 110 147
rect 113 145 115 147
rect 185 145 187 147
rect 190 145 192 147
rect 195 145 197 147
rect 200 145 202 147
rect 205 145 207 147
rect 210 145 212 147
rect 215 145 217 147
rect 220 145 222 147
rect 225 145 227 147
rect 230 145 232 147
rect 235 145 237 147
rect 240 145 242 147
rect 248 145 250 147
rect 253 145 255 147
rect 258 145 260 147
rect 273 144 275 146
rect 20 139 22 141
rect 40 140 42 142
rect 45 140 47 142
rect 50 140 52 142
rect 248 140 250 142
rect 253 140 255 142
rect 258 140 260 142
rect 273 139 275 141
rect 20 134 22 136
rect 40 135 42 137
rect 45 135 47 137
rect 50 135 52 137
rect 248 135 250 137
rect 253 135 255 137
rect 258 135 260 137
rect 273 134 275 136
rect 20 129 22 131
rect 40 130 42 132
rect 45 130 47 132
rect 50 130 52 132
rect 248 130 250 132
rect 253 130 255 132
rect 258 130 260 132
rect 273 129 275 131
rect 146 127 148 129
rect 151 127 153 129
rect 20 124 22 126
rect 40 125 42 127
rect 45 125 47 127
rect 50 125 52 127
rect 248 125 250 127
rect 253 125 255 127
rect 258 125 260 127
rect 273 124 275 126
rect 20 119 22 121
rect 40 120 42 122
rect 45 120 47 122
rect 50 120 52 122
rect 248 120 250 122
rect 253 120 255 122
rect 258 120 260 122
rect 273 119 275 121
rect 20 114 22 116
rect 40 115 42 117
rect 45 115 47 117
rect 50 115 52 117
rect 248 115 250 117
rect 253 115 255 117
rect 258 115 260 117
rect 273 114 275 116
rect 20 109 22 111
rect 40 110 42 112
rect 45 110 47 112
rect 50 110 52 112
rect 58 110 60 112
rect 63 110 65 112
rect 68 110 70 112
rect 73 110 75 112
rect 78 110 80 112
rect 83 110 85 112
rect 88 110 90 112
rect 93 110 95 112
rect 98 110 100 112
rect 103 110 105 112
rect 108 110 110 112
rect 113 110 115 112
rect 185 110 187 112
rect 190 110 192 112
rect 195 110 197 112
rect 200 110 202 112
rect 205 110 207 112
rect 210 110 212 112
rect 215 110 217 112
rect 220 110 222 112
rect 225 110 227 112
rect 230 110 232 112
rect 235 110 237 112
rect 240 110 242 112
rect 248 110 250 112
rect 253 110 255 112
rect 258 110 260 112
rect 273 109 275 111
rect 20 104 22 106
rect 273 104 275 106
rect 20 99 22 101
rect 273 99 275 101
rect 20 94 22 96
rect 273 94 275 96
rect 20 89 22 91
rect 273 89 275 91
rect 20 84 22 86
rect 273 84 275 86
rect 20 79 22 81
rect 40 80 42 82
rect 45 80 47 82
rect 50 80 52 82
rect 58 80 60 82
rect 63 80 65 82
rect 68 80 70 82
rect 73 80 75 82
rect 78 80 80 82
rect 83 80 85 82
rect 88 80 90 82
rect 93 80 95 82
rect 98 80 100 82
rect 103 80 105 82
rect 108 80 110 82
rect 113 80 115 82
rect 185 80 187 82
rect 190 80 192 82
rect 195 80 197 82
rect 200 80 202 82
rect 205 80 207 82
rect 210 80 212 82
rect 215 80 217 82
rect 220 80 222 82
rect 225 80 227 82
rect 230 80 232 82
rect 235 80 237 82
rect 240 80 242 82
rect 248 80 250 82
rect 253 80 255 82
rect 258 80 260 82
rect 273 79 275 81
rect 20 74 22 76
rect 40 75 42 77
rect 45 75 47 77
rect 50 75 52 77
rect 248 75 250 77
rect 253 75 255 77
rect 258 75 260 77
rect 273 74 275 76
rect 20 69 22 71
rect 40 70 42 72
rect 45 70 47 72
rect 50 70 52 72
rect 248 70 250 72
rect 253 70 255 72
rect 258 70 260 72
rect 273 69 275 71
rect 20 64 22 66
rect 40 65 42 67
rect 45 65 47 67
rect 50 65 52 67
rect 248 65 250 67
rect 253 65 255 67
rect 258 65 260 67
rect 146 63 148 65
rect 151 63 153 65
rect 273 64 275 66
rect 20 59 22 61
rect 40 60 42 62
rect 45 60 47 62
rect 50 60 52 62
rect 248 60 250 62
rect 253 60 255 62
rect 258 60 260 62
rect 273 59 275 61
rect 20 54 22 56
rect 40 55 42 57
rect 45 55 47 57
rect 50 55 52 57
rect 146 55 148 57
rect 151 55 153 57
rect 248 55 250 57
rect 253 55 255 57
rect 258 55 260 57
rect 273 54 275 56
rect 20 49 22 51
rect 40 50 42 52
rect 45 50 47 52
rect 50 50 52 52
rect 248 50 250 52
rect 253 50 255 52
rect 258 50 260 52
rect 273 49 275 51
rect 146 47 148 49
rect 151 47 153 49
rect 20 44 22 46
rect 40 45 42 47
rect 45 45 47 47
rect 50 45 52 47
rect 58 45 60 47
rect 63 45 65 47
rect 68 45 70 47
rect 73 45 75 47
rect 78 45 80 47
rect 83 45 85 47
rect 88 45 90 47
rect 93 45 95 47
rect 205 45 207 47
rect 210 45 212 47
rect 215 45 217 47
rect 220 45 222 47
rect 225 45 227 47
rect 230 45 232 47
rect 235 45 237 47
rect 240 45 242 47
rect 248 45 250 47
rect 253 45 255 47
rect 258 45 260 47
rect 273 44 275 46
rect 20 39 22 41
rect 146 39 148 41
rect 151 39 153 41
rect 273 39 275 41
rect 20 34 22 36
rect 273 34 275 36
rect 146 31 148 33
rect 151 31 153 33
rect 20 29 22 31
rect 40 29 42 31
rect 45 29 47 31
rect 50 29 52 31
rect 55 29 57 31
rect 60 29 62 31
rect 65 29 67 31
rect 70 29 72 31
rect 75 29 77 31
rect 80 29 82 31
rect 85 29 87 31
rect 90 29 92 31
rect 95 29 97 31
rect 203 29 205 31
rect 208 29 210 31
rect 213 29 215 31
rect 218 29 220 31
rect 223 29 225 31
rect 228 29 230 31
rect 233 29 235 31
rect 238 29 240 31
rect 243 29 245 31
rect 248 29 250 31
rect 253 29 255 31
rect 258 29 260 31
rect 273 29 275 31
rect 20 18 22 20
rect 25 18 27 20
rect 30 18 32 20
rect 35 18 37 20
rect 40 18 42 20
rect 45 18 47 20
rect 50 18 52 20
rect 55 18 57 20
rect 60 18 62 20
rect 65 18 67 20
rect 70 18 72 20
rect 75 18 77 20
rect 80 18 82 20
rect 85 18 87 20
rect 90 18 92 20
rect 95 18 97 20
rect 203 18 205 20
rect 208 18 210 20
rect 213 18 215 20
rect 218 18 220 20
rect 223 18 225 20
rect 228 18 230 20
rect 233 18 235 20
rect 238 18 240 20
rect 243 18 245 20
rect 248 18 250 20
rect 253 18 255 20
rect 258 18 260 20
rect 263 18 265 20
rect 268 18 270 20
rect 273 18 275 20
rect 278 18 280 20
<< metal3 >>
rect 23 743 277 997
<< gv2 >>
rect 47 971 49 973
rect 59 971 61 973
rect 71 971 73 973
rect 83 971 85 973
rect 95 971 97 973
rect 107 971 109 973
rect 119 971 121 973
rect 131 971 133 973
rect 143 971 145 973
rect 155 971 157 973
rect 167 971 169 973
rect 179 971 181 973
rect 191 971 193 973
rect 203 971 205 973
rect 215 971 217 973
rect 227 971 229 973
rect 239 971 241 973
rect 251 971 253 973
rect 47 959 49 961
rect 59 959 61 961
rect 71 959 73 961
rect 83 959 85 961
rect 95 959 97 961
rect 107 959 109 961
rect 119 959 121 961
rect 131 959 133 961
rect 143 959 145 961
rect 155 959 157 961
rect 167 959 169 961
rect 179 959 181 961
rect 191 959 193 961
rect 203 959 205 961
rect 215 959 217 961
rect 227 959 229 961
rect 239 959 241 961
rect 251 959 253 961
rect 47 947 49 949
rect 59 947 61 949
rect 71 947 73 949
rect 83 947 85 949
rect 95 947 97 949
rect 107 947 109 949
rect 119 947 121 949
rect 131 947 133 949
rect 143 947 145 949
rect 155 947 157 949
rect 167 947 169 949
rect 179 947 181 949
rect 191 947 193 949
rect 203 947 205 949
rect 215 947 217 949
rect 227 947 229 949
rect 239 947 241 949
rect 251 947 253 949
rect 47 935 49 937
rect 59 935 61 937
rect 71 935 73 937
rect 83 935 85 937
rect 95 935 97 937
rect 107 935 109 937
rect 119 935 121 937
rect 131 935 133 937
rect 143 935 145 937
rect 155 935 157 937
rect 167 935 169 937
rect 179 935 181 937
rect 191 935 193 937
rect 203 935 205 937
rect 215 935 217 937
rect 227 935 229 937
rect 239 935 241 937
rect 251 935 253 937
rect 47 923 49 925
rect 59 923 61 925
rect 71 923 73 925
rect 83 923 85 925
rect 95 923 97 925
rect 107 923 109 925
rect 119 923 121 925
rect 131 923 133 925
rect 143 923 145 925
rect 155 923 157 925
rect 167 923 169 925
rect 179 923 181 925
rect 191 923 193 925
rect 203 923 205 925
rect 215 923 217 925
rect 227 923 229 925
rect 239 923 241 925
rect 251 923 253 925
rect 47 911 49 913
rect 59 911 61 913
rect 71 911 73 913
rect 83 911 85 913
rect 95 911 97 913
rect 107 911 109 913
rect 119 911 121 913
rect 131 911 133 913
rect 143 911 145 913
rect 155 911 157 913
rect 167 911 169 913
rect 179 911 181 913
rect 191 911 193 913
rect 203 911 205 913
rect 215 911 217 913
rect 227 911 229 913
rect 239 911 241 913
rect 251 911 253 913
rect 47 899 49 901
rect 59 899 61 901
rect 71 899 73 901
rect 83 899 85 901
rect 95 899 97 901
rect 107 899 109 901
rect 119 899 121 901
rect 131 899 133 901
rect 143 899 145 901
rect 155 899 157 901
rect 167 899 169 901
rect 179 899 181 901
rect 191 899 193 901
rect 203 899 205 901
rect 215 899 217 901
rect 227 899 229 901
rect 239 899 241 901
rect 251 899 253 901
rect 47 887 49 889
rect 59 887 61 889
rect 71 887 73 889
rect 83 887 85 889
rect 95 887 97 889
rect 107 887 109 889
rect 119 887 121 889
rect 131 887 133 889
rect 143 887 145 889
rect 155 887 157 889
rect 167 887 169 889
rect 179 887 181 889
rect 191 887 193 889
rect 203 887 205 889
rect 215 887 217 889
rect 227 887 229 889
rect 239 887 241 889
rect 251 887 253 889
rect 47 875 49 877
rect 59 875 61 877
rect 71 875 73 877
rect 83 875 85 877
rect 95 875 97 877
rect 107 875 109 877
rect 119 875 121 877
rect 131 875 133 877
rect 143 875 145 877
rect 155 875 157 877
rect 167 875 169 877
rect 179 875 181 877
rect 191 875 193 877
rect 203 875 205 877
rect 215 875 217 877
rect 227 875 229 877
rect 239 875 241 877
rect 251 875 253 877
rect 47 863 49 865
rect 59 863 61 865
rect 71 863 73 865
rect 83 863 85 865
rect 95 863 97 865
rect 107 863 109 865
rect 119 863 121 865
rect 131 863 133 865
rect 143 863 145 865
rect 155 863 157 865
rect 167 863 169 865
rect 179 863 181 865
rect 191 863 193 865
rect 203 863 205 865
rect 215 863 217 865
rect 227 863 229 865
rect 239 863 241 865
rect 251 863 253 865
rect 47 851 49 853
rect 59 851 61 853
rect 71 851 73 853
rect 83 851 85 853
rect 95 851 97 853
rect 107 851 109 853
rect 119 851 121 853
rect 131 851 133 853
rect 143 851 145 853
rect 155 851 157 853
rect 167 851 169 853
rect 179 851 181 853
rect 191 851 193 853
rect 203 851 205 853
rect 215 851 217 853
rect 227 851 229 853
rect 239 851 241 853
rect 251 851 253 853
rect 47 839 49 841
rect 59 839 61 841
rect 71 839 73 841
rect 83 839 85 841
rect 95 839 97 841
rect 107 839 109 841
rect 119 839 121 841
rect 131 839 133 841
rect 143 839 145 841
rect 155 839 157 841
rect 167 839 169 841
rect 179 839 181 841
rect 191 839 193 841
rect 203 839 205 841
rect 215 839 217 841
rect 227 839 229 841
rect 239 839 241 841
rect 251 839 253 841
rect 47 827 49 829
rect 59 827 61 829
rect 71 827 73 829
rect 83 827 85 829
rect 95 827 97 829
rect 107 827 109 829
rect 119 827 121 829
rect 131 827 133 829
rect 143 827 145 829
rect 155 827 157 829
rect 167 827 169 829
rect 179 827 181 829
rect 191 827 193 829
rect 203 827 205 829
rect 215 827 217 829
rect 227 827 229 829
rect 239 827 241 829
rect 251 827 253 829
rect 47 815 49 817
rect 59 815 61 817
rect 71 815 73 817
rect 83 815 85 817
rect 95 815 97 817
rect 107 815 109 817
rect 119 815 121 817
rect 131 815 133 817
rect 143 815 145 817
rect 155 815 157 817
rect 167 815 169 817
rect 179 815 181 817
rect 191 815 193 817
rect 203 815 205 817
rect 215 815 217 817
rect 227 815 229 817
rect 239 815 241 817
rect 251 815 253 817
rect 47 803 49 805
rect 59 803 61 805
rect 71 803 73 805
rect 83 803 85 805
rect 95 803 97 805
rect 107 803 109 805
rect 119 803 121 805
rect 131 803 133 805
rect 143 803 145 805
rect 155 803 157 805
rect 167 803 169 805
rect 179 803 181 805
rect 191 803 193 805
rect 203 803 205 805
rect 215 803 217 805
rect 227 803 229 805
rect 239 803 241 805
rect 251 803 253 805
rect 47 791 49 793
rect 59 791 61 793
rect 71 791 73 793
rect 83 791 85 793
rect 95 791 97 793
rect 107 791 109 793
rect 119 791 121 793
rect 131 791 133 793
rect 143 791 145 793
rect 155 791 157 793
rect 167 791 169 793
rect 179 791 181 793
rect 191 791 193 793
rect 203 791 205 793
rect 215 791 217 793
rect 227 791 229 793
rect 239 791 241 793
rect 251 791 253 793
rect 47 779 49 781
rect 59 779 61 781
rect 71 779 73 781
rect 83 779 85 781
rect 95 779 97 781
rect 107 779 109 781
rect 119 779 121 781
rect 131 779 133 781
rect 143 779 145 781
rect 155 779 157 781
rect 167 779 169 781
rect 179 779 181 781
rect 191 779 193 781
rect 203 779 205 781
rect 215 779 217 781
rect 227 779 229 781
rect 239 779 241 781
rect 251 779 253 781
rect 47 767 49 769
rect 59 767 61 769
rect 71 767 73 769
rect 83 767 85 769
rect 95 767 97 769
rect 107 767 109 769
rect 119 767 121 769
rect 131 767 133 769
rect 143 767 145 769
rect 155 767 157 769
rect 167 767 169 769
rect 179 767 181 769
rect 191 767 193 769
rect 203 767 205 769
rect 215 767 217 769
rect 227 767 229 769
rect 239 767 241 769
rect 251 767 253 769
<< glass >>
rect 43 763 257 977
<< xp >>
rect 23 743 277 997
<< labels >>
rlabel metal1 150 -1 150 -1 8 Vdd!
rlabel metal2 140 126 140 126 6 gnd:2
rlabel metal1 150 -9 150 -9 8 Vdd!
<< end >>
