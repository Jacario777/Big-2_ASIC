magic
tech scmos
timestamp 1681620392
<< metal1 >>
rect -762 4730 -701 4765
rect -457 4725 -404 4764
rect -160 4723 -105 4767
rect 136 4725 201 4762
rect 438 4730 501 4765
rect 738 4728 806 4764
rect 1037 4726 1102 4758
rect 1342 4729 1399 4766
rect 1635 4732 1710 4763
rect 1938 4726 2001 4764
rect 2244 4729 2300 4759
rect 2541 4723 2597 4769
rect 2837 4725 2901 4761
rect 3136 4722 3202 4764
rect 3438 4724 3502 4763
rect 3739 4726 3798 4767
rect -858 4016 -852 4019
rect -858 4015 -846 4016
rect -858 4013 -844 4015
rect -858 4010 -839 4013
rect -558 4010 -552 4019
rect -258 4010 -252 4019
rect 42 4010 48 4019
rect 1021 4010 1117 4026
rect 1542 4010 1548 4019
rect 1842 4010 1848 4019
rect 2142 4010 2148 4019
rect 2442 4010 2448 4019
rect 2742 4010 2748 4019
rect 3126 4018 3212 4026
rect 3131 4010 3207 4018
rect 3342 4010 3348 4019
rect 3642 4010 3648 4019
rect -858 4007 3889 4010
rect -855 4006 3889 4007
rect -853 4004 3889 4006
rect -851 4001 3889 4004
rect -851 3995 1112 4001
rect -1610 3853 -1572 3916
rect -851 3767 -839 3995
rect 1026 3993 1112 3995
rect 342 3980 348 3986
rect 642 3980 648 3986
rect 1031 3985 1107 3993
rect 3141 3992 3889 4001
rect -862 3761 -839 3767
rect -1610 3553 -1574 3619
rect -1614 3314 -1577 3321
rect -1614 3253 -1573 3314
rect -1614 3252 -1577 3253
rect -1612 2961 -1567 3013
rect -851 2816 -839 3761
rect -823 3962 960 3980
rect 1036 3977 1102 3985
rect 1242 3980 1248 3986
rect 1041 3969 1097 3977
rect -823 3467 -805 3962
rect -829 3461 -805 3467
rect -823 3167 -805 3461
rect -829 3161 -805 3167
rect -823 2867 -805 3161
rect 1046 3027 1092 3969
rect 1178 3962 3058 3980
rect 3141 3326 3197 3992
rect 3271 3962 3855 3980
rect 2547 3270 3197 3326
rect 2547 3027 2603 3270
rect 14 3007 3077 3027
rect 38 2983 3053 3003
rect 38 2967 3053 2973
rect -829 2861 -805 2867
rect -870 2726 -862 2731
rect -1608 2661 -1564 2722
rect -870 2721 -854 2726
rect -870 2716 -846 2721
rect -870 2710 -838 2716
rect -823 2710 -805 2861
rect -134 2901 58 2946
rect 426 2943 452 2946
rect 426 2936 429 2943
rect 1610 2936 1613 2945
rect 364 2933 372 2936
rect 386 2926 389 2935
rect 412 2933 429 2936
rect 466 2933 508 2936
rect 148 2923 173 2926
rect 204 2923 221 2926
rect 324 2923 341 2926
rect 380 2923 389 2926
rect 466 2925 469 2933
rect 554 2926 557 2935
rect 610 2933 628 2936
rect 692 2933 717 2936
rect 796 2933 821 2936
rect 836 2933 861 2936
rect 882 2926 885 2935
rect 986 2933 996 2936
rect 1010 2933 1020 2936
rect 1058 2926 1061 2935
rect 1178 2933 1188 2936
rect 1202 2926 1205 2935
rect 1522 2926 1525 2935
rect 1538 2933 1548 2936
rect 1572 2933 1581 2936
rect 1610 2933 1628 2936
rect 1642 2933 1660 2936
rect 2010 2933 2028 2936
rect 2154 2926 2157 2935
rect 2170 2933 2180 2936
rect 2204 2933 2213 2936
rect 2226 2926 2229 2935
rect 2754 2926 2757 2935
rect 2882 2933 2892 2936
rect 538 2923 557 2926
rect 676 2923 684 2926
rect 802 2923 828 2926
rect 834 2923 876 2926
rect 882 2923 892 2926
rect 1004 2923 1021 2926
rect 1036 2923 1052 2926
rect 1058 2923 1068 2926
rect 1162 2923 1172 2926
rect 1196 2923 1205 2926
rect 1266 2923 1276 2926
rect 1452 2923 1477 2926
rect 1508 2923 1525 2926
rect 1532 2923 1549 2926
rect 1570 2923 1588 2926
rect 1636 2923 1661 2926
rect 1722 2923 1748 2926
rect 1948 2923 1973 2926
rect 2026 2923 2036 2926
rect 2148 2923 2157 2926
rect 2202 2923 2220 2926
rect 2226 2923 2236 2926
rect 2266 2923 2292 2926
rect 2372 2923 2381 2926
rect 2692 2923 2701 2926
rect 2748 2923 2757 2926
rect 2874 2923 2900 2926
rect 228 2913 237 2916
rect 284 2913 317 2916
rect 338 2915 341 2923
rect 698 2913 724 2916
rect 1018 2915 1021 2923
rect 1546 2915 1549 2923
rect 2202 2915 2205 2923
rect 258 2903 276 2906
rect -134 2710 -89 2901
rect 3033 2895 3198 2940
rect 14 2867 3077 2873
rect 114 2833 140 2836
rect 258 2833 276 2836
rect 780 2833 797 2836
rect 260 2823 269 2826
rect 284 2823 317 2826
rect 522 2823 540 2826
rect 844 2823 853 2826
rect 1132 2823 1141 2826
rect 1252 2823 1261 2826
rect 1324 2823 1333 2826
rect 850 2816 853 2823
rect 1594 2816 1597 2825
rect 1914 2816 1917 2825
rect 1988 2823 1997 2826
rect 1994 2816 1997 2823
rect 2050 2816 2053 2825
rect 2226 2816 2229 2825
rect 2378 2816 2381 2825
rect 2834 2816 2837 2825
rect 356 2813 373 2816
rect 378 2806 381 2814
rect 466 2813 484 2816
rect 516 2813 533 2816
rect 562 2813 573 2816
rect 642 2813 660 2816
rect 692 2813 709 2816
rect 850 2813 876 2816
rect 882 2813 900 2816
rect 1076 2813 1109 2816
rect 1138 2813 1148 2816
rect 1218 2813 1236 2816
rect 1250 2813 1284 2816
rect 1290 2813 1308 2816
rect 1356 2813 1365 2816
rect 1444 2813 1469 2816
rect 1500 2813 1509 2816
rect 1516 2813 1525 2816
rect 1564 2813 1573 2816
rect 1580 2813 1597 2816
rect 1636 2813 1661 2816
rect 1682 2813 1700 2816
rect 1706 2813 1724 2816
rect 1858 2813 1876 2816
rect 1914 2813 1932 2816
rect 1994 2813 2012 2816
rect 2050 2813 2068 2816
rect 2074 2813 2092 2816
rect 2122 2813 2148 2816
rect 2226 2813 2244 2816
rect 2250 2813 2260 2816
rect 2290 2813 2316 2816
rect 2378 2813 2396 2816
rect 2410 2813 2428 2816
rect 2452 2813 2469 2816
rect 2546 2813 2572 2816
rect 2586 2813 2596 2816
rect 2602 2813 2620 2816
rect 2788 2813 2797 2816
rect 2820 2813 2837 2816
rect 2908 2813 2917 2816
rect 466 2806 469 2813
rect 202 2803 228 2806
rect 322 2803 332 2806
rect 364 2803 381 2806
rect 410 2803 420 2806
rect 452 2803 469 2806
rect 492 2803 501 2806
rect 570 2805 573 2813
rect 596 2803 613 2806
rect 634 2803 668 2806
rect 706 2805 709 2813
rect 748 2803 765 2806
rect 882 2805 885 2813
rect 994 2803 1004 2806
rect 1018 2803 1028 2806
rect 1178 2803 1196 2806
rect 1218 2805 1221 2813
rect 1252 2803 1269 2806
rect 1362 2805 1365 2813
rect 1506 2805 1509 2813
rect 1538 2803 1556 2806
rect 1562 2803 1572 2806
rect 1642 2803 1660 2806
rect 1684 2803 1693 2806
rect 1826 2803 1836 2806
rect 1882 2803 1892 2806
rect 1938 2803 1964 2806
rect 2052 2803 2061 2806
rect 2074 2805 2077 2813
rect 2194 2803 2204 2806
rect 2228 2803 2237 2806
rect 2250 2805 2253 2813
rect 2404 2803 2421 2806
rect 2458 2803 2468 2806
rect 2492 2803 2501 2806
rect 2546 2805 2549 2813
rect 2554 2803 2564 2806
rect 2794 2805 2797 2813
rect 2860 2803 2869 2806
rect 290 2793 324 2796
rect 1530 2793 1548 2796
rect 38 2767 3053 2773
rect 164 2743 173 2746
rect 1266 2743 1284 2746
rect 146 2733 156 2736
rect 180 2733 189 2736
rect 338 2733 348 2736
rect 396 2733 405 2736
rect 474 2733 500 2736
rect 524 2733 533 2736
rect 570 2733 580 2736
rect 602 2726 605 2735
rect 610 2733 628 2736
rect 794 2726 797 2735
rect 810 2733 820 2736
rect 1164 2733 1189 2736
rect 1212 2733 1236 2736
rect 1300 2733 1324 2736
rect 1516 2733 1533 2736
rect 242 2723 252 2726
rect 356 2723 365 2726
rect 482 2723 508 2726
rect 522 2723 548 2726
rect 564 2723 581 2726
rect 602 2723 613 2726
rect 634 2723 652 2726
rect 732 2723 757 2726
rect 788 2723 797 2726
rect 804 2723 821 2726
rect 836 2723 845 2726
rect 866 2723 876 2726
rect 996 2723 1005 2726
rect 1172 2723 1181 2726
rect 1186 2725 1189 2733
rect 1658 2726 1661 2735
rect 2018 2726 2021 2735
rect 2346 2726 2349 2735
rect 2892 2733 2901 2736
rect 1220 2723 1228 2726
rect 1308 2723 1316 2726
rect 1340 2723 1357 2726
rect 1428 2723 1453 2726
rect 1508 2723 1548 2726
rect 1652 2723 1661 2726
rect 1860 2723 1885 2726
rect 2012 2723 2021 2726
rect 2164 2723 2173 2726
rect 2260 2723 2285 2726
rect 2346 2723 2364 2726
rect 2834 2723 2844 2726
rect 2866 2723 2876 2726
rect 2890 2723 2908 2726
rect 468 2713 493 2716
rect 818 2715 821 2723
rect 1354 2715 1357 2723
rect 2890 2715 2893 2723
rect -870 2665 -89 2710
rect 442 2703 460 2706
rect 1682 2703 1692 2706
rect 1714 2703 1724 2706
rect 1770 2703 1788 2706
rect 14 2667 3077 2673
rect -870 2660 -838 2665
rect -870 2655 -846 2660
rect -870 2650 -854 2655
rect -870 2645 -862 2650
rect -851 2515 -839 2558
rect -862 2509 -839 2515
rect -1610 2359 -1566 2416
rect -1606 2066 -1571 2111
rect -851 1967 -839 2509
rect -862 1961 -839 1967
rect -1615 1765 -1571 1814
rect -851 1667 -839 1961
rect -862 1661 -839 1667
rect -1606 1455 -1570 1520
rect -1605 1162 -1564 1212
rect -851 1025 -839 1661
rect -823 1367 -811 2665
rect 546 2633 564 2636
rect 548 2623 557 2626
rect 572 2623 581 2626
rect 842 2616 845 2625
rect 1170 2616 1173 2625
rect 1260 2623 1269 2626
rect 1346 2623 1364 2626
rect 1498 2616 1501 2625
rect 2730 2623 2764 2626
rect 2866 2616 2869 2625
rect 108 2613 133 2616
rect 164 2613 173 2616
rect 292 2613 309 2616
rect 346 2613 356 2616
rect 370 2613 412 2616
rect 468 2613 477 2616
rect 586 2613 596 2616
rect 828 2613 845 2616
rect 988 2613 1005 2616
rect 1044 2613 1069 2616
rect 1100 2613 1109 2616
rect 1170 2613 1181 2616
rect 1202 2613 1212 2616
rect 1218 2613 1244 2616
rect 1266 2613 1284 2616
rect 1306 2613 1324 2616
rect 1354 2613 1372 2616
rect 1378 2613 1396 2616
rect 1410 2613 1428 2616
rect 1484 2613 1501 2616
rect 1516 2613 1541 2616
rect 1786 2613 1796 2616
rect 1868 2613 1877 2616
rect 2042 2613 2060 2616
rect 2114 2613 2124 2616
rect 2186 2613 2196 2616
rect 2202 2613 2244 2616
rect 2258 2613 2269 2616
rect 2276 2613 2285 2616
rect 2324 2613 2332 2616
rect 2370 2613 2380 2616
rect 2434 2613 2444 2616
rect 2532 2613 2541 2616
rect 2786 2613 2852 2616
rect 2866 2613 2884 2616
rect 170 2605 173 2613
rect 260 2603 268 2606
rect 364 2603 405 2606
rect 490 2603 500 2606
rect 684 2603 701 2606
rect 834 2603 844 2606
rect 1106 2605 1109 2613
rect 1132 2603 1141 2606
rect 1178 2605 1181 2613
rect 1220 2603 1229 2606
rect 1490 2603 1500 2606
rect 2042 2605 2045 2613
rect 2068 2603 2077 2606
rect 372 2593 381 2596
rect 666 2593 676 2596
rect 2114 2593 2117 2613
rect 2122 2603 2132 2606
rect 2148 2603 2157 2606
rect 2186 2605 2189 2613
rect 2204 2603 2221 2606
rect 2226 2603 2236 2606
rect 2266 2605 2269 2613
rect 2356 2603 2372 2606
rect 2436 2603 2445 2606
rect 2468 2603 2484 2606
rect 2594 2603 2604 2606
rect 2660 2603 2677 2606
rect 2786 2605 2789 2613
rect 2868 2603 2877 2606
rect 2892 2603 2917 2606
rect 38 2567 3053 2573
rect 1012 2543 1020 2546
rect 170 2526 173 2534
rect 108 2523 133 2526
rect 164 2523 173 2526
rect 180 2523 189 2526
rect 234 2523 237 2534
rect 250 2523 253 2534
rect 282 2526 285 2534
rect 418 2526 421 2534
rect 658 2533 676 2536
rect 978 2533 1004 2536
rect 1018 2533 1028 2536
rect 1050 2526 1053 2534
rect 1140 2533 1157 2536
rect 1162 2533 1172 2536
rect 1202 2533 1212 2536
rect 1226 2533 1236 2536
rect 1378 2533 1404 2536
rect 1546 2526 1549 2534
rect 1962 2533 1972 2536
rect 2018 2533 2028 2536
rect 2044 2533 2053 2536
rect 2132 2533 2148 2536
rect 2644 2533 2653 2536
rect 2700 2533 2717 2536
rect 2892 2533 2901 2536
rect 258 2523 276 2526
rect 282 2523 308 2526
rect 402 2523 412 2526
rect 418 2523 428 2526
rect 474 2523 484 2526
rect 522 2523 532 2526
rect 692 2523 709 2526
rect 810 2523 820 2526
rect 1044 2523 1053 2526
rect 1060 2523 1077 2526
rect 1090 2523 1116 2526
rect 1220 2523 1229 2526
rect 1260 2523 1269 2526
rect 1420 2523 1445 2526
rect 1476 2523 1493 2526
rect 1508 2523 1549 2526
rect 1690 2523 1700 2526
rect 1714 2523 1732 2526
rect 1850 2523 1860 2526
rect 1874 2523 1884 2526
rect 2002 2523 2020 2526
rect 2060 2523 2077 2526
rect 2092 2523 2101 2526
rect 2202 2523 2220 2526
rect 2268 2523 2277 2526
rect 2316 2523 2325 2526
rect 2612 2523 2621 2526
rect 2658 2523 2676 2526
rect 2850 2523 2876 2526
rect 2890 2523 2908 2526
rect 652 2513 661 2516
rect 666 2513 676 2516
rect 1434 2513 1468 2516
rect 1490 2515 1493 2523
rect 2714 2513 2724 2516
rect 2890 2515 2893 2523
rect 3153 2509 3198 2895
rect 3837 2509 3855 3962
rect 3871 3767 3889 3992
rect 4601 3859 4646 3911
rect 3871 3761 3900 3767
rect 3871 3467 3889 3761
rect 4601 3564 4643 3611
rect 3871 3461 3900 3467
rect 3871 3167 3889 3461
rect 4603 3259 4648 3312
rect 3871 3161 3900 3167
rect 3871 2867 3889 3161
rect 4602 2968 4649 3011
rect 3871 2861 3900 2867
rect 3871 2567 3889 2861
rect 4610 2669 4644 2715
rect 3871 2561 3900 2567
rect 3871 2552 3889 2561
rect 842 2503 868 2506
rect 14 2467 3077 2473
rect 3153 2464 3860 2509
rect 212 2433 252 2436
rect 442 2433 460 2436
rect 722 2433 748 2436
rect 228 2423 236 2426
rect 434 2423 453 2426
rect 468 2423 485 2426
rect 722 2423 732 2426
rect 756 2423 764 2426
rect 836 2423 844 2426
rect 932 2423 941 2426
rect 434 2416 437 2423
rect 1602 2416 1605 2425
rect 1866 2423 1876 2426
rect 2202 2416 2205 2425
rect 2330 2423 2340 2426
rect 2410 2423 2436 2426
rect 2498 2423 2532 2426
rect 2562 2423 2572 2426
rect 2674 2423 2716 2426
rect 2330 2416 2333 2423
rect 2410 2416 2413 2423
rect 2826 2416 2829 2425
rect 2850 2423 2900 2426
rect 66 2413 76 2416
rect 66 2403 69 2413
rect 242 2403 245 2414
rect 308 2413 317 2416
rect 338 2413 356 2416
rect 362 2413 372 2416
rect 428 2413 437 2416
rect 586 2413 596 2416
rect 602 2413 628 2416
rect 786 2413 828 2416
rect 972 2413 989 2416
rect 996 2413 1012 2416
rect 1026 2413 1036 2416
rect 1060 2413 1077 2416
rect 1124 2413 1149 2416
rect 1180 2413 1197 2416
rect 1204 2413 1213 2416
rect 1372 2413 1381 2416
rect 1468 2413 1493 2416
rect 1540 2413 1557 2416
rect 1578 2413 1588 2416
rect 1602 2413 1620 2416
rect 1802 2413 1812 2416
rect 1836 2413 1845 2416
rect 1860 2413 1877 2416
rect 2036 2413 2053 2416
rect 2114 2413 2140 2416
rect 2202 2413 2220 2416
rect 2250 2413 2260 2416
rect 2308 2413 2333 2416
rect 2356 2413 2365 2416
rect 2396 2413 2413 2416
rect 2476 2413 2517 2416
rect 2562 2413 2580 2416
rect 2602 2413 2636 2416
rect 276 2403 285 2406
rect 380 2403 389 2406
rect 396 2403 405 2406
rect 420 2403 429 2406
rect 604 2403 613 2406
rect 938 2403 964 2406
rect 978 2403 988 2406
rect 1010 2403 1020 2406
rect 1194 2405 1197 2413
rect 2690 2406 2693 2416
rect 2738 2413 2756 2416
rect 2778 2413 2812 2416
rect 2826 2413 2844 2416
rect 2874 2413 2908 2416
rect 3815 2411 3860 2464
rect 3900 2426 3908 2431
rect 3892 2421 3908 2426
rect 3884 2416 3908 2421
rect 3876 2411 3908 2416
rect 1236 2403 1260 2406
rect 1546 2403 1556 2406
rect 1570 2403 1580 2406
rect 1844 2403 1853 2406
rect 2042 2403 2052 2406
rect 2226 2403 2236 2406
rect 2282 2403 2300 2406
rect 2322 2403 2340 2406
rect 2364 2403 2373 2406
rect 2484 2403 2525 2406
rect 2556 2403 2573 2406
rect 2594 2403 2628 2406
rect 2676 2403 2693 2406
rect 2706 2403 2716 2406
rect 2852 2403 2885 2406
rect 386 2395 389 2403
rect 1242 2393 1252 2396
rect 38 2367 3053 2373
rect 3815 2366 3908 2411
rect 3876 2360 3908 2366
rect 3884 2355 3908 2360
rect 4605 2356 4646 2422
rect 3892 2350 3908 2355
rect 66 2343 84 2346
rect 3900 2345 3908 2350
rect 66 2333 92 2336
rect 156 2333 165 2336
rect 108 2323 117 2326
rect 124 2323 133 2326
rect 274 2325 277 2336
rect 186 2313 196 2316
rect 210 2313 220 2316
rect 226 2306 229 2315
rect 234 2313 237 2325
rect 290 2323 300 2326
rect 322 2323 340 2326
rect 386 2325 389 2336
rect 402 2323 405 2334
rect 444 2333 452 2336
rect 684 2333 693 2336
rect 876 2333 893 2336
rect 1050 2326 1053 2334
rect 1292 2333 1301 2336
rect 1564 2333 1572 2336
rect 2394 2326 2397 2334
rect 2442 2326 2445 2334
rect 2482 2333 2524 2336
rect 436 2323 453 2326
rect 564 2323 573 2326
rect 682 2323 692 2326
rect 804 2323 813 2326
rect 818 2323 844 2326
rect 860 2323 869 2326
rect 1012 2323 1029 2326
rect 1050 2323 1068 2326
rect 1074 2323 1092 2326
rect 1234 2323 1252 2326
rect 1258 2323 1284 2326
rect 1370 2323 1380 2326
rect 1436 2323 1445 2326
rect 1618 2323 1644 2326
rect 1756 2323 1765 2326
rect 1836 2323 1844 2326
rect 1924 2323 1933 2326
rect 2020 2323 2045 2326
rect 2116 2323 2141 2326
rect 2220 2323 2237 2326
rect 2372 2323 2397 2326
rect 2404 2323 2429 2326
rect 2434 2323 2445 2326
rect 2452 2323 2461 2326
rect 2476 2323 2501 2326
rect 2540 2323 2549 2326
rect 2564 2323 2573 2326
rect 2588 2323 2597 2326
rect 2636 2323 2661 2326
rect 348 2313 357 2316
rect 420 2313 428 2316
rect 468 2313 485 2316
rect 538 2313 548 2316
rect 924 2313 933 2316
rect 1018 2313 1028 2316
rect 1682 2313 1700 2316
rect 204 2303 229 2306
rect 482 2306 485 2313
rect 482 2303 508 2306
rect 890 2303 916 2306
rect 14 2267 3077 2273
rect 842 2233 861 2236
rect 474 2223 484 2226
rect 842 2216 845 2233
rect 66 2213 76 2216
rect 122 2213 132 2216
rect 212 2213 237 2216
rect 268 2213 277 2216
rect 284 2213 293 2216
rect 274 2205 277 2213
rect 314 2206 317 2216
rect 362 2206 365 2216
rect 500 2213 516 2216
rect 562 2213 588 2216
rect 644 2213 660 2216
rect 314 2205 325 2206
rect 316 2203 325 2205
rect 362 2203 372 2206
rect 810 2205 813 2216
rect 836 2213 845 2216
rect 858 2215 861 2233
rect 1090 2226 1093 2236
rect 1298 2233 1332 2236
rect 876 2223 885 2226
rect 972 2223 981 2226
rect 1084 2223 1093 2226
rect 1138 2216 1141 2225
rect 1242 2223 1260 2226
rect 1274 2223 1284 2226
rect 1450 2223 1460 2226
rect 1562 2223 1572 2226
rect 1594 2216 1597 2225
rect 1740 2223 1748 2226
rect 2090 2216 2093 2225
rect 2122 2216 2125 2225
rect 2146 2216 2149 2225
rect 2234 2216 2237 2225
rect 2314 2216 2317 2225
rect 2596 2223 2604 2226
rect 2698 2216 2701 2225
rect 2948 2223 2965 2226
rect 2970 2223 2980 2226
rect 2962 2216 2965 2223
rect 906 2213 916 2216
rect 940 2213 949 2216
rect 964 2213 973 2216
rect 1004 2213 1013 2216
rect 882 2203 892 2206
rect 922 2203 932 2206
rect 946 2203 956 2206
rect 1044 2203 1053 2206
rect 1090 2205 1093 2216
rect 1100 2213 1117 2216
rect 1138 2213 1148 2216
rect 1220 2213 1229 2216
rect 1236 2213 1253 2216
rect 1370 2213 1381 2216
rect 1444 2213 1461 2216
rect 1468 2213 1485 2216
rect 1492 2213 1501 2216
rect 1580 2213 1597 2216
rect 1716 2213 1725 2216
rect 1804 2213 1821 2216
rect 1884 2213 1892 2216
rect 1980 2213 1989 2216
rect 2090 2213 2108 2216
rect 2114 2213 2125 2216
rect 2132 2213 2149 2216
rect 2188 2213 2205 2216
rect 2234 2213 2252 2216
rect 2258 2213 2277 2216
rect 2282 2213 2300 2216
rect 2314 2213 2332 2216
rect 2476 2213 2485 2216
rect 2538 2213 2548 2216
rect 2554 2213 2581 2216
rect 2612 2213 2645 2216
rect 2698 2213 2716 2216
rect 2764 2213 2781 2216
rect 2962 2213 2988 2216
rect 1106 2203 1116 2206
rect 1378 2205 1381 2213
rect 1722 2205 1725 2213
rect 2258 2205 2261 2213
rect 2266 2203 2292 2206
rect 2554 2205 2557 2213
rect 2562 2203 2580 2206
rect 2620 2203 2629 2206
rect 2642 2203 2660 2206
rect 2666 2203 2676 2206
rect 2948 2203 2957 2206
rect 2996 2203 3013 2206
rect 1026 2193 1036 2196
rect 38 2167 3053 2173
rect 802 2143 820 2146
rect 220 2133 229 2136
rect 700 2133 725 2136
rect 788 2133 821 2136
rect 828 2133 845 2136
rect 898 2133 908 2136
rect 954 2133 964 2136
rect 978 2133 988 2136
rect 1154 2133 1172 2136
rect 1228 2133 1237 2136
rect 1244 2133 1261 2136
rect 108 2123 125 2126
rect 180 2123 189 2126
rect 266 2123 292 2126
rect 364 2123 389 2126
rect 444 2123 460 2126
rect 522 2123 540 2126
rect 612 2123 629 2126
rect 698 2123 732 2126
rect 738 2123 756 2126
rect 762 2123 772 2126
rect 892 2123 909 2126
rect 916 2123 925 2126
rect 972 2123 981 2126
rect 1274 2125 1277 2136
rect 1626 2126 1629 2135
rect 1658 2133 1668 2136
rect 1692 2133 1717 2136
rect 2196 2133 2213 2136
rect 2348 2133 2381 2136
rect 2404 2133 2437 2136
rect 2682 2133 2692 2136
rect 2714 2133 2724 2136
rect 2738 2133 2756 2136
rect 2802 2133 2812 2136
rect 2836 2133 2845 2136
rect 1316 2123 1333 2126
rect 1428 2123 1453 2126
rect 1564 2123 1589 2126
rect 1620 2123 1629 2126
rect 1780 2123 1804 2126
rect 1818 2123 1836 2126
rect 1884 2123 1909 2126
rect 1940 2123 1949 2126
rect 1970 2123 1988 2126
rect 2060 2123 2085 2126
rect 2116 2123 2125 2126
rect 2322 2123 2332 2126
rect 2378 2123 2396 2126
rect 2444 2123 2461 2126
rect 2482 2123 2500 2126
rect 2514 2123 2524 2126
rect 2716 2123 2725 2126
rect 2732 2123 2757 2126
rect 2778 2123 2796 2126
rect 2834 2123 2852 2126
rect 2988 2123 2997 2126
rect 700 2113 709 2116
rect 788 2113 813 2116
rect 924 2113 965 2116
rect 980 2113 989 2116
rect 1268 2113 1277 2116
rect 1292 2113 1300 2116
rect 1818 2115 1821 2123
rect 1970 2115 1973 2123
rect 2378 2116 2381 2123
rect 1996 2113 2004 2116
rect 2196 2113 2205 2116
rect 2348 2113 2381 2116
rect 2410 2113 2436 2116
rect 2482 2115 2485 2123
rect 2778 2115 2781 2123
rect 2834 2115 2837 2123
rect 1186 2103 1204 2106
rect 1266 2103 1284 2106
rect 14 2067 3077 2073
rect 522 2016 525 2025
rect 1234 2023 1244 2026
rect 1618 2016 1621 2025
rect 2498 2023 2508 2026
rect 2682 2016 2685 2025
rect 2988 2023 2996 2026
rect 66 2013 76 2016
rect 138 2013 148 2016
rect 154 2013 180 2016
rect 236 2013 261 2016
rect 266 2013 276 2016
rect 522 2013 532 2016
rect 538 2013 565 2016
rect 612 2013 637 2016
rect 138 2005 141 2013
rect 826 2006 829 2014
rect 156 2003 165 2006
rect 204 2003 237 2006
rect 242 2003 268 2006
rect 490 2003 500 2006
rect 764 2003 829 2006
rect 858 2006 861 2014
rect 858 2003 884 2006
rect 890 2003 893 2014
rect 924 2013 957 2016
rect 1252 2013 1285 2016
rect 1322 2013 1348 2016
rect 1436 2013 1461 2016
rect 1492 2013 1501 2016
rect 1596 2013 1621 2016
rect 1684 2013 1709 2016
rect 1818 2013 1844 2016
rect 1916 2013 1933 2016
rect 1972 2013 1981 2016
rect 2042 2013 2076 2016
rect 2132 2013 2157 2016
rect 2188 2013 2197 2016
rect 2244 2013 2269 2016
rect 2300 2013 2309 2016
rect 2316 2013 2325 2016
rect 2396 2013 2421 2016
rect 2506 2013 2516 2016
rect 2676 2013 2685 2016
rect 2700 2013 2709 2016
rect 898 2003 908 2006
rect 922 2003 956 2006
rect 1212 2003 1245 2006
rect 1498 2005 1501 2013
rect 1580 2003 1588 2006
rect 1602 2003 1620 2006
rect 1978 2005 1981 2013
rect 1994 2003 2012 2006
rect 2058 2003 2068 2006
rect 2194 2005 2197 2013
rect 2306 2005 2309 2013
rect 2322 2005 2325 2013
rect 2524 2003 2549 2006
rect 2650 2003 2668 2006
rect 2708 2003 2717 2006
rect 2786 2003 2796 2006
rect 2802 2003 2805 2014
rect 2812 2013 2829 2016
rect 2842 2013 2852 2016
rect 2908 2013 2917 2016
rect 2970 2013 2980 2016
rect 2994 2013 3004 2016
rect 234 1996 237 2003
rect 234 1993 261 1996
rect 866 1993 876 1996
rect 924 1993 933 1996
rect 38 1967 3053 1973
rect 3871 1967 3889 2253
rect 4605 2066 4647 2111
rect 3871 1961 3900 1967
rect 234 1943 268 1946
rect 82 1933 100 1936
rect 130 1933 156 1936
rect 210 1926 213 1935
rect 234 1933 276 1936
rect 354 1933 364 1936
rect 492 1933 501 1936
rect 562 1933 572 1936
rect 82 1923 92 1926
rect 130 1923 148 1926
rect 180 1923 189 1926
rect 194 1923 204 1926
rect 210 1923 221 1926
rect 234 1925 237 1933
rect 602 1926 605 1935
rect 858 1926 861 1935
rect 970 1933 980 1936
rect 1082 1933 1092 1936
rect 1490 1926 1493 1935
rect 1524 1933 1572 1936
rect 2010 1926 2013 1935
rect 2026 1926 2029 1935
rect 2260 1933 2293 1936
rect 2434 1926 2437 1935
rect 2450 1933 2476 1936
rect 2524 1933 2541 1936
rect 2666 1933 2676 1936
rect 2700 1933 2709 1936
rect 2730 1933 2756 1936
rect 356 1923 372 1926
rect 508 1923 517 1926
rect 596 1923 605 1926
rect 852 1923 861 1926
rect 956 1923 973 1926
rect 1004 1923 1045 1926
rect 1082 1923 1109 1926
rect 1162 1923 1172 1926
rect 1306 1923 1332 1926
rect 1412 1923 1437 1926
rect 1468 1923 1493 1926
rect 1500 1923 1509 1926
rect 1516 1923 1525 1926
rect 1588 1923 1605 1926
rect 1644 1923 1668 1926
rect 1708 1923 1733 1926
rect 1810 1923 1820 1926
rect 1834 1923 1852 1926
rect 1858 1923 1892 1926
rect 2010 1923 2020 1926
rect 2026 1923 2036 1926
rect 2066 1923 2092 1926
rect 2156 1923 2165 1926
rect 2236 1923 2285 1926
rect 2428 1923 2437 1926
rect 2474 1923 2484 1926
rect 2498 1923 2509 1926
rect 2516 1923 2533 1926
rect 2692 1923 2701 1926
rect 2764 1923 2773 1926
rect 2786 1923 2796 1926
rect 404 1913 412 1916
rect 490 1913 500 1916
rect 1018 1913 1052 1916
rect 1082 1906 1085 1923
rect 1122 1913 1132 1916
rect 1530 1913 1572 1916
rect 1834 1915 1837 1923
rect 1860 1913 1869 1916
rect 2498 1915 2501 1923
rect 378 1903 396 1906
rect 882 1903 892 1906
rect 1060 1903 1085 1906
rect 1252 1903 1269 1906
rect 14 1867 3077 1873
rect 908 1833 925 1836
rect 1122 1833 1132 1836
rect 372 1823 381 1826
rect 890 1823 900 1826
rect 914 1823 933 1826
rect 1450 1816 1453 1825
rect 1546 1816 1549 1825
rect 2602 1823 2612 1826
rect 2794 1823 2804 1826
rect 2868 1823 2885 1826
rect 2882 1816 2885 1823
rect 2914 1816 2917 1825
rect 106 1813 116 1816
rect 122 1813 156 1816
rect 196 1813 204 1816
rect 226 1813 236 1816
rect 242 1813 260 1816
rect 308 1813 325 1816
rect 340 1813 364 1816
rect 442 1813 460 1816
rect 474 1813 492 1816
rect 564 1813 581 1816
rect 756 1813 765 1816
rect 812 1813 837 1816
rect 868 1813 877 1816
rect 884 1813 893 1816
rect 1004 1813 1013 1816
rect 1050 1813 1076 1816
rect 1146 1813 1156 1816
rect 1306 1813 1316 1816
rect 1370 1813 1388 1816
rect 1394 1813 1404 1816
rect 124 1803 141 1806
rect 212 1803 228 1806
rect 314 1803 324 1806
rect 498 1803 516 1806
rect 972 1803 980 1806
rect 1340 1803 1349 1806
rect 1362 1803 1380 1806
rect 1426 1805 1429 1816
rect 1450 1813 1468 1816
rect 1522 1813 1532 1816
rect 1538 1813 1549 1816
rect 1634 1813 1652 1816
rect 1868 1813 1877 1816
rect 1900 1813 1917 1816
rect 1948 1813 1964 1816
rect 2020 1813 2029 1816
rect 2116 1813 2141 1816
rect 2172 1813 2181 1816
rect 1540 1803 1549 1806
rect 1722 1803 1740 1806
rect 1874 1805 1877 1813
rect 1906 1803 1924 1806
rect 1972 1803 1989 1806
rect 2178 1805 2181 1813
rect 2330 1805 2333 1816
rect 2364 1813 2373 1816
rect 2468 1813 2477 1816
rect 2490 1813 2500 1816
rect 2474 1805 2477 1813
rect 2506 1805 2509 1816
rect 2626 1813 2636 1816
rect 2532 1803 2541 1806
rect 2588 1803 2605 1806
rect 2626 1805 2629 1813
rect 2658 1806 2661 1814
rect 2666 1813 2676 1816
rect 2690 1813 2701 1816
rect 2658 1803 2668 1806
rect 2690 1805 2693 1813
rect 2714 1805 2717 1816
rect 2724 1813 2741 1816
rect 2730 1803 2748 1806
rect 2770 1805 2773 1816
rect 2810 1805 2813 1816
rect 2842 1805 2845 1816
rect 2866 1805 2869 1816
rect 2882 1813 2908 1816
rect 2914 1813 2932 1816
rect 2874 1803 2900 1806
rect 2914 1803 2924 1806
rect 2948 1803 2957 1806
rect 38 1767 3053 1773
rect 658 1743 684 1746
rect 698 1743 708 1746
rect 722 1743 732 1746
rect 1170 1743 1180 1746
rect 1236 1743 1244 1746
rect 314 1733 324 1736
rect 386 1726 389 1735
rect 426 1733 452 1736
rect 546 1733 564 1736
rect 426 1726 429 1733
rect 546 1726 549 1733
rect 188 1723 205 1726
rect 386 1723 397 1726
rect 412 1723 429 1726
rect 434 1723 460 1726
rect 522 1723 549 1726
rect 594 1726 597 1735
rect 618 1733 644 1736
rect 692 1733 701 1736
rect 716 1733 733 1736
rect 594 1723 685 1726
rect 700 1723 709 1726
rect 748 1723 765 1726
rect 812 1723 821 1726
rect 826 1716 829 1735
rect 842 1733 852 1736
rect 890 1733 900 1736
rect 1052 1733 1060 1736
rect 890 1725 893 1733
rect 1098 1726 1101 1735
rect 1188 1733 1197 1736
rect 1228 1733 1245 1736
rect 1252 1733 1284 1736
rect 1410 1733 1420 1736
rect 1586 1726 1589 1735
rect 1604 1733 1620 1736
rect 1634 1733 1644 1736
rect 1666 1733 1676 1736
rect 1700 1733 1741 1736
rect 1778 1726 1781 1735
rect 1834 1733 1844 1736
rect 2258 1726 2261 1735
rect 2282 1733 2308 1736
rect 2340 1733 2373 1736
rect 2754 1733 2764 1736
rect 2810 1733 2852 1736
rect 2898 1726 2901 1735
rect 956 1723 973 1726
rect 1012 1723 1021 1726
rect 1084 1723 1101 1726
rect 1146 1723 1164 1726
rect 1204 1723 1220 1726
rect 1322 1723 1332 1726
rect 1338 1723 1349 1726
rect 1396 1723 1405 1726
rect 1428 1723 1453 1726
rect 1586 1723 1596 1726
rect 1628 1723 1645 1726
rect 1652 1723 1661 1726
rect 1666 1723 1684 1726
rect 1778 1723 1845 1726
rect 1866 1723 1884 1726
rect 1932 1723 1941 1726
rect 2100 1723 2125 1726
rect 2252 1723 2261 1726
rect 2268 1723 2277 1726
rect 2332 1723 2349 1726
rect 2532 1723 2557 1726
rect 2618 1723 2636 1726
rect 2804 1723 2813 1726
rect 2860 1723 2869 1726
rect 2874 1723 2884 1726
rect 2898 1723 2909 1726
rect 354 1713 364 1716
rect 820 1713 829 1716
rect 1346 1716 1349 1723
rect 1346 1713 1356 1716
rect 1700 1713 1733 1716
rect 1346 1703 1372 1706
rect 14 1667 3077 1673
rect 3871 1667 3889 1961
rect 4608 1765 4647 1814
rect 3871 1661 3900 1667
rect 1570 1633 1580 1636
rect 1650 1633 1668 1636
rect 2828 1633 2845 1636
rect 938 1623 948 1626
rect 108 1613 133 1616
rect 244 1613 253 1616
rect 250 1606 253 1613
rect 330 1613 340 1616
rect 346 1613 356 1616
rect 386 1613 412 1616
rect 484 1613 501 1616
rect 578 1613 596 1616
rect 602 1613 612 1616
rect 666 1613 709 1616
rect 204 1603 213 1606
rect 250 1603 260 1606
rect 330 1605 333 1613
rect 346 1605 349 1613
rect 578 1605 581 1613
rect 620 1603 637 1606
rect 644 1603 677 1606
rect 706 1605 709 1613
rect 722 1603 725 1614
rect 748 1613 781 1616
rect 788 1613 829 1616
rect 892 1613 901 1616
rect 1020 1613 1037 1616
rect 1114 1613 1132 1616
rect 754 1603 780 1606
rect 802 1603 828 1606
rect 1114 1605 1117 1613
rect 1234 1606 1237 1625
rect 1148 1603 1165 1606
rect 1172 1603 1189 1606
rect 1204 1603 1237 1606
rect 1258 1603 1276 1606
rect 1290 1603 1293 1625
rect 1300 1623 1309 1626
rect 1506 1623 1516 1626
rect 1676 1623 1684 1626
rect 2604 1623 2613 1626
rect 2730 1616 2733 1625
rect 2844 1623 2853 1626
rect 1330 1613 1340 1616
rect 1442 1613 1460 1616
rect 1532 1613 1549 1616
rect 1620 1613 1629 1616
rect 1692 1613 1701 1616
rect 1740 1613 1765 1616
rect 1964 1613 1972 1616
rect 2140 1613 2165 1616
rect 2196 1613 2213 1616
rect 2276 1613 2301 1616
rect 2332 1613 2341 1616
rect 2508 1613 2517 1616
rect 2540 1613 2548 1616
rect 2602 1613 2620 1616
rect 2634 1613 2668 1616
rect 2698 1613 2716 1616
rect 2730 1613 2748 1616
rect 1386 1603 1404 1606
rect 1546 1605 1549 1613
rect 2068 1603 2077 1606
rect 2098 1603 2116 1606
rect 2338 1605 2341 1613
rect 2506 1603 2524 1606
rect 2604 1603 2612 1606
rect 2684 1603 2701 1606
rect 2834 1603 2837 1614
rect 2874 1613 2884 1616
rect 2890 1613 2908 1616
rect 628 1593 636 1596
rect 1156 1593 1164 1596
rect 38 1567 3053 1573
rect 290 1543 300 1546
rect 314 1543 340 1546
rect 1082 1543 1108 1546
rect 1122 1543 1132 1546
rect 186 1526 189 1534
rect 242 1533 284 1536
rect 378 1533 412 1536
rect 538 1533 556 1536
rect 108 1523 133 1526
rect 178 1523 189 1526
rect 236 1523 269 1526
rect 292 1523 301 1526
rect 316 1523 341 1526
rect 386 1523 404 1526
rect 418 1523 436 1526
rect 466 1523 492 1526
rect 570 1525 573 1536
rect 580 1533 613 1536
rect 636 1533 693 1536
rect 714 1533 724 1536
rect 762 1533 772 1536
rect 802 1533 836 1536
rect 850 1533 860 1536
rect 882 1533 900 1536
rect 986 1533 1012 1536
rect 1068 1533 1077 1536
rect 586 1523 628 1526
rect 690 1515 693 1533
rect 1082 1526 1085 1543
rect 1116 1533 1133 1536
rect 1140 1533 1196 1536
rect 1210 1533 1220 1536
rect 1260 1533 1292 1536
rect 1386 1533 1412 1536
rect 1538 1533 1564 1536
rect 1578 1526 1581 1534
rect 2178 1526 2181 1534
rect 2244 1533 2253 1536
rect 2268 1533 2277 1536
rect 2450 1533 2484 1536
rect 2602 1533 2621 1536
rect 2626 1526 2629 1534
rect 2820 1533 2837 1536
rect 700 1523 709 1526
rect 740 1523 765 1526
rect 770 1523 780 1526
rect 844 1523 861 1526
rect 868 1523 893 1526
rect 970 1523 980 1526
rect 986 1523 1020 1526
rect 1042 1523 1085 1526
rect 1124 1523 1133 1526
rect 1204 1523 1221 1526
rect 1252 1523 1277 1526
rect 1306 1523 1317 1526
rect 1324 1523 1333 1526
rect 1386 1523 1404 1526
rect 1506 1523 1565 1526
rect 1572 1523 1581 1526
rect 1618 1523 1628 1526
rect 1658 1523 1684 1526
rect 1732 1523 1748 1526
rect 1802 1523 1828 1526
rect 2020 1523 2037 1526
rect 2116 1523 2133 1526
rect 2172 1523 2181 1526
rect 2210 1523 2228 1526
rect 2242 1523 2260 1526
rect 2396 1523 2420 1526
rect 2434 1523 2444 1526
rect 2482 1523 2492 1526
rect 2618 1523 2629 1526
rect 2748 1523 2764 1526
rect 2804 1523 2812 1526
rect 2914 1523 2948 1526
rect 788 1513 837 1516
rect 930 1513 940 1516
rect 1236 1513 1244 1516
rect 1306 1515 1309 1523
rect 1330 1516 1333 1523
rect 1330 1513 1356 1516
rect 1434 1513 1452 1516
rect 1482 1513 1516 1516
rect 2242 1515 2245 1523
rect 2866 1513 2876 1516
rect 938 1503 956 1506
rect 14 1467 3077 1473
rect 418 1433 444 1436
rect 1266 1433 1292 1436
rect 218 1423 228 1426
rect 242 1423 276 1426
rect 290 1423 300 1426
rect 452 1423 509 1426
rect 524 1423 533 1426
rect 858 1416 861 1425
rect 890 1423 916 1426
rect 1010 1416 1013 1425
rect 1266 1416 1269 1433
rect 1386 1423 1420 1426
rect 2124 1423 2141 1426
rect 156 1413 165 1416
rect 202 1413 236 1416
rect 274 1413 284 1416
rect 308 1413 333 1416
rect 340 1413 357 1416
rect 364 1413 397 1416
rect 516 1413 541 1416
rect 618 1413 644 1416
rect 90 1403 148 1406
rect 162 1405 165 1413
rect 188 1403 229 1406
rect 244 1403 253 1406
rect 498 1403 508 1406
rect 522 1403 548 1406
rect 722 1405 725 1416
rect 738 1413 764 1416
rect 788 1413 813 1416
rect 820 1413 837 1416
rect 858 1413 868 1416
rect 956 1413 988 1416
rect 1002 1413 1013 1416
rect 1076 1413 1101 1416
rect 1138 1413 1148 1416
rect 1252 1413 1269 1416
rect 1428 1413 1453 1416
rect 1468 1413 1477 1416
rect 1554 1413 1580 1416
rect 1820 1413 1845 1416
rect 1876 1413 1885 1416
rect 1892 1413 1940 1416
rect 2052 1413 2069 1416
rect 2130 1413 2180 1416
rect 802 1403 812 1406
rect 834 1405 837 1413
rect 970 1403 980 1406
rect 1002 1405 1005 1413
rect 1172 1403 1189 1406
rect 1380 1403 1389 1406
rect 1436 1403 1460 1406
rect 1474 1403 1484 1406
rect 1882 1405 1885 1413
rect 1906 1403 1932 1406
rect 2082 1403 2092 1406
rect 2122 1403 2172 1406
rect 2202 1405 2205 1416
rect 2252 1413 2277 1416
rect 2332 1413 2397 1416
rect 2418 1406 2421 1425
rect 2452 1423 2461 1426
rect 2860 1423 2885 1426
rect 2882 1416 2885 1423
rect 2484 1413 2493 1416
rect 2500 1413 2517 1416
rect 2546 1413 2556 1416
rect 2418 1403 2428 1406
rect 2458 1403 2476 1406
rect 2578 1405 2581 1416
rect 2666 1413 2676 1416
rect 2724 1413 2733 1416
rect 2764 1413 2781 1416
rect 2786 1413 2796 1416
rect 2882 1413 2916 1416
rect 2922 1413 2932 1416
rect 2938 1406 2941 1425
rect 2962 1423 2972 1426
rect 2988 1413 3005 1416
rect 2770 1403 2788 1406
rect 2860 1403 2869 1406
rect 2874 1403 2908 1406
rect 2938 1403 2972 1406
rect 38 1367 3053 1373
rect 3871 1367 3889 1661
rect 4609 1460 4649 1519
rect -829 1361 -811 1367
rect -823 1067 -811 1361
rect 3871 1361 3900 1367
rect 108 1343 125 1346
rect 2874 1343 2908 1346
rect 122 1326 125 1343
rect 162 1333 173 1336
rect 250 1333 276 1336
rect 324 1333 340 1336
rect 122 1323 132 1326
rect 162 1325 165 1333
rect 530 1326 533 1334
rect 690 1326 693 1334
rect 186 1323 220 1326
rect 258 1323 284 1326
rect 322 1323 332 1326
rect 370 1323 380 1326
rect 442 1323 452 1326
rect 492 1323 501 1326
rect 516 1323 533 1326
rect 554 1323 564 1326
rect 684 1323 693 1326
rect 770 1325 773 1336
rect 794 1323 797 1334
rect 804 1323 829 1326
rect 850 1325 853 1336
rect 194 1313 212 1316
rect 298 1313 308 1316
rect 554 1315 557 1323
rect 826 1313 836 1316
rect 410 1303 428 1306
rect 826 1293 829 1313
rect 866 1306 869 1334
rect 882 1333 924 1336
rect 938 1333 956 1336
rect 994 1333 1004 1336
rect 1172 1333 1188 1336
rect 1226 1326 1229 1334
rect 1252 1333 1269 1336
rect 1292 1333 1301 1336
rect 1402 1333 1428 1336
rect 1450 1326 1453 1334
rect 1476 1333 1485 1336
rect 1634 1326 1637 1334
rect 1818 1326 1821 1334
rect 876 1323 925 1326
rect 932 1323 949 1326
rect 1148 1323 1156 1326
rect 1218 1323 1229 1326
rect 1244 1323 1284 1326
rect 1436 1323 1453 1326
rect 1474 1323 1500 1326
rect 1628 1323 1637 1326
rect 1660 1323 1676 1326
rect 1708 1323 1717 1326
rect 1756 1323 1781 1326
rect 1812 1323 1821 1326
rect 1908 1323 1925 1326
rect 1964 1323 1973 1326
rect 2028 1323 2053 1326
rect 2090 1323 2093 1334
rect 2124 1333 2132 1336
rect 2162 1323 2165 1334
rect 2266 1326 2269 1334
rect 2386 1326 2389 1334
rect 2260 1323 2269 1326
rect 2380 1323 2389 1326
rect 2458 1323 2461 1334
rect 2642 1323 2645 1334
rect 2810 1333 2836 1336
rect 2916 1333 2932 1336
rect 2946 1333 2988 1336
rect 2746 1323 2764 1326
rect 2796 1323 2821 1326
rect 2834 1323 2844 1326
rect 2930 1323 2940 1326
rect 2996 1323 3005 1326
rect 1218 1316 1221 1323
rect 1212 1313 1221 1316
rect 1290 1313 1316 1316
rect 1340 1313 1349 1316
rect 1692 1313 1700 1316
rect 2818 1313 2821 1323
rect 844 1303 869 1306
rect 1298 1303 1332 1306
rect 14 1267 3077 1273
rect 106 1233 140 1236
rect 234 1233 253 1236
rect 114 1223 124 1226
rect 114 1216 117 1223
rect 92 1213 117 1216
rect 234 1215 237 1233
rect 250 1225 253 1233
rect 418 1233 461 1236
rect 1348 1233 1365 1236
rect 1644 1233 1653 1236
rect 340 1223 349 1226
rect 324 1213 333 1216
rect 370 1213 380 1216
rect 418 1215 421 1233
rect 458 1215 461 1233
rect 476 1223 493 1226
rect 578 1216 581 1225
rect 1330 1223 1340 1226
rect 1674 1223 1684 1226
rect 2322 1216 2325 1225
rect 500 1213 525 1216
rect 540 1213 549 1216
rect 170 1203 188 1206
rect 482 1203 492 1206
rect 522 1203 525 1213
rect 546 1205 549 1213
rect 570 1213 581 1216
rect 740 1213 765 1216
rect 796 1213 805 1216
rect 812 1213 828 1216
rect 570 1205 573 1213
rect 802 1205 805 1213
rect 882 1205 885 1216
rect 980 1213 989 1216
rect 1092 1213 1101 1216
rect 1196 1213 1221 1216
rect 1252 1213 1261 1216
rect 1282 1213 1300 1216
rect 986 1205 989 1213
rect 1098 1205 1101 1213
rect 1148 1203 1157 1206
rect 1258 1205 1261 1213
rect 1324 1203 1333 1206
rect 1410 1205 1413 1216
rect 1548 1213 1573 1216
rect 1762 1213 1788 1216
rect 1826 1213 1836 1216
rect 1898 1213 1916 1216
rect 1620 1203 1629 1206
rect 1930 1205 1933 1216
rect 2068 1213 2093 1216
rect 2124 1213 2133 1216
rect 2140 1213 2156 1216
rect 2268 1213 2277 1216
rect 2314 1213 2325 1216
rect 2130 1205 2133 1213
rect 2346 1205 2349 1216
rect 2354 1205 2357 1216
rect 2412 1213 2437 1216
rect 2498 1205 2501 1216
rect 2610 1213 2620 1216
rect 2634 1213 2652 1216
rect 2682 1213 2732 1216
rect 2762 1213 2772 1216
rect 2812 1214 2820 1216
rect 2810 1213 2820 1214
rect 2852 1213 2885 1216
rect 2668 1203 2693 1206
rect 2706 1203 2724 1206
rect 2788 1203 2797 1206
rect 2810 1203 2813 1213
rect 2882 1206 2885 1213
rect 2818 1203 2828 1206
rect 2866 1205 2885 1206
rect 2866 1203 2884 1205
rect 38 1167 3053 1173
rect 250 1143 276 1146
rect 290 1143 300 1146
rect 1524 1143 1533 1146
rect 1674 1136 1677 1145
rect 284 1133 301 1136
rect 338 1133 380 1136
rect 554 1126 557 1135
rect 818 1133 844 1136
rect 860 1133 869 1136
rect 874 1133 892 1136
rect 1034 1126 1037 1135
rect 1516 1133 1533 1136
rect 1650 1133 1660 1136
rect 1674 1133 1684 1136
rect 1530 1126 1533 1133
rect 1714 1126 1717 1135
rect 1740 1133 1765 1136
rect 1866 1126 1869 1135
rect 1898 1126 1901 1136
rect 1922 1133 1932 1136
rect 1956 1133 1965 1136
rect 1980 1133 1997 1136
rect 2658 1133 2676 1136
rect 2698 1133 2732 1136
rect 2754 1133 2796 1136
rect 2890 1133 2900 1136
rect 2922 1133 2932 1136
rect 2946 1133 2972 1136
rect 108 1123 133 1126
rect 164 1123 181 1126
rect 228 1123 237 1126
rect 332 1123 373 1126
rect 404 1123 413 1126
rect 450 1123 476 1126
rect 546 1123 557 1126
rect 572 1123 613 1126
rect 674 1123 700 1126
rect 826 1123 836 1126
rect 868 1123 884 1126
rect 972 1123 997 1126
rect 1028 1123 1037 1126
rect 1116 1123 1141 1126
rect 1362 1123 1372 1126
rect 1436 1123 1477 1126
rect 1530 1123 1548 1126
rect 1554 1123 1588 1126
rect 1618 1123 1652 1126
rect 1692 1123 1717 1126
rect 1804 1123 1829 1126
rect 1860 1123 1869 1126
rect 1876 1123 1940 1126
rect 1954 1123 1972 1126
rect 2036 1123 2061 1126
rect 2124 1123 2148 1126
rect 2266 1123 2276 1126
rect 2434 1123 2444 1126
rect 2794 1123 2804 1126
rect 2940 1123 2965 1126
rect 2988 1123 3005 1126
rect 170 1113 188 1116
rect 642 1113 652 1116
rect 1380 1113 1397 1116
rect 1402 1113 1428 1116
rect 1740 1113 1749 1116
rect 1954 1115 1957 1123
rect 2962 1116 2965 1123
rect 2962 1113 2972 1116
rect 14 1067 3077 1073
rect 3871 1067 3889 1361
rect 4605 1156 4650 1214
rect -829 1061 -811 1067
rect -870 926 -862 931
rect -870 921 -854 926
rect -1607 852 -1564 920
rect -870 916 -846 921
rect -870 910 -838 916
rect -823 910 -811 1061
rect 3871 1061 3900 1067
rect 426 1033 436 1036
rect 482 1033 500 1036
rect 444 1023 453 1026
rect 1668 1023 1677 1026
rect 1692 1023 1701 1026
rect 1884 1023 1909 1026
rect 2188 1023 2197 1026
rect 2386 1023 2404 1026
rect 2884 1023 2893 1026
rect 2940 1023 2949 1026
rect 210 1013 228 1016
rect 276 1013 309 1016
rect 314 1006 317 1014
rect 356 1013 373 1016
rect 380 1013 389 1016
rect 404 1013 413 1016
rect 186 1003 220 1006
rect 244 1003 261 1006
rect 274 1003 317 1006
rect 364 1003 372 1006
rect 722 1005 725 1016
rect 738 1013 756 1016
rect 762 1013 813 1016
rect 860 1013 869 1016
rect 890 1013 900 1016
rect 938 1013 964 1016
rect 1058 1013 1084 1016
rect 1098 1013 1108 1016
rect 1148 1013 1157 1016
rect 780 1003 805 1006
rect 818 1003 836 1006
rect 858 1003 868 1006
rect 930 1003 956 1006
rect 986 1003 1028 1006
rect 1100 1003 1109 1006
rect 1132 1003 1141 1006
rect 1156 1003 1165 1006
rect 1276 1003 1293 1006
rect 1330 1003 1333 1014
rect 1444 1013 1461 1016
rect 1516 1013 1525 1016
rect 1684 1013 1693 1016
rect 1458 1005 1461 1013
rect 1514 1003 1556 1006
rect 1642 1003 1652 1006
rect 1666 1003 1676 1006
rect 1698 1005 1701 1023
rect 2386 1016 2389 1023
rect 1730 1003 1733 1014
rect 1804 1013 1813 1016
rect 1866 1005 1869 1016
rect 1876 1013 1901 1016
rect 1948 1013 1973 1016
rect 2004 1013 2021 1016
rect 2028 1013 2044 1016
rect 2090 1013 2109 1016
rect 2116 1013 2125 1016
rect 2132 1013 2141 1016
rect 2146 1013 2172 1016
rect 2292 1013 2301 1016
rect 2332 1013 2349 1016
rect 2356 1013 2389 1016
rect 2420 1013 2461 1016
rect 2562 1013 2580 1016
rect 2620 1013 2645 1016
rect 2018 1005 2021 1013
rect 2068 1003 2101 1006
rect 2106 1005 2109 1013
rect 2154 1003 2164 1006
rect 2188 1003 2197 1006
rect 2338 1003 2348 1006
rect 2394 1003 2404 1006
rect 2428 1003 2437 1006
rect 2634 1003 2652 1006
rect 2674 1005 2677 1016
rect 2682 1005 2685 1016
rect 2692 1013 2709 1016
rect 2730 1013 2748 1016
rect 2698 1003 2708 1006
rect 2770 1005 2773 1016
rect 2804 1013 2853 1016
rect 2906 1013 2924 1016
rect 2812 1003 2837 1006
rect 2850 1003 2860 1006
rect 2970 1003 2988 1006
rect 250 993 260 996
rect 38 967 3053 973
rect 218 943 236 946
rect 2996 943 3013 946
rect 204 933 213 936
rect 244 933 277 936
rect 322 926 325 935
rect 412 933 420 936
rect 1082 926 1085 935
rect 1098 933 1116 936
rect 1202 926 1205 935
rect 1274 933 1308 936
rect 1330 926 1333 936
rect 1364 933 1389 936
rect 1418 933 1436 936
rect 1458 933 1492 936
rect 1522 933 1540 936
rect 1554 933 1564 936
rect 1578 933 1596 936
rect 1610 933 1620 936
rect 1634 935 1644 936
rect 1634 933 1645 935
rect 1642 926 1645 933
rect 108 923 133 926
rect 292 923 325 926
rect 332 923 341 926
rect 356 923 365 926
rect 386 923 397 926
rect 404 923 421 926
rect 428 923 445 926
rect 602 923 612 926
rect 692 923 701 926
rect 772 923 781 926
rect 972 923 981 926
rect 1076 923 1085 926
rect 1106 923 1124 926
rect 1164 923 1205 926
rect 1242 923 1268 926
rect 1330 925 1349 926
rect 1332 923 1349 925
rect 1362 923 1388 926
rect 1460 923 1484 926
rect 1548 923 1565 926
rect 1572 923 1597 926
rect 1604 923 1621 926
rect 1628 923 1645 926
rect 1666 926 1669 935
rect 1690 926 1693 935
rect 1756 933 1773 936
rect 1826 926 1829 935
rect 1844 933 1861 936
rect 1866 933 1876 936
rect 2180 933 2189 936
rect 2324 933 2348 936
rect 2386 933 2396 936
rect 2418 926 2421 935
rect 2436 933 2477 936
rect 2610 926 2613 935
rect 2626 933 2636 936
rect 2674 933 2708 936
rect 2988 933 3005 936
rect 1666 923 1677 926
rect 1684 923 1693 926
rect 1722 923 1740 926
rect 1826 923 1877 926
rect 2052 923 2077 926
rect 2140 923 2164 926
rect 2178 923 2196 926
rect 2356 923 2397 926
rect 2418 923 2469 926
rect 2604 923 2613 926
rect 2620 923 2644 926
rect 2860 923 2877 926
rect 2938 923 2956 926
rect 2962 923 2980 926
rect 300 913 317 916
rect 394 915 397 923
rect 442 916 445 923
rect 1242 916 1245 923
rect 442 913 452 916
rect 476 913 485 916
rect 540 913 549 916
rect 652 913 661 916
rect 940 913 949 916
rect 1228 913 1245 916
rect 1276 913 1293 916
rect 1762 913 1772 916
rect 2178 915 2181 923
rect 2378 913 2396 916
rect 2442 913 2484 916
rect 2898 913 2908 916
rect 2938 915 2941 923
rect -870 865 -99 910
rect 442 903 468 906
rect 538 903 556 906
rect 650 903 668 906
rect 14 867 3077 873
rect -870 860 -838 865
rect -870 855 -846 860
rect -870 850 -854 855
rect -870 845 -862 850
rect -1607 560 -1569 613
rect -1606 268 -1565 308
rect -851 167 -839 761
rect -862 161 -839 167
rect -1608 -42 -1568 19
rect -851 -30 -839 161
rect -823 -3 -805 865
rect -144 436 -99 865
rect 2914 833 2932 836
rect 380 823 389 826
rect 522 823 548 826
rect 850 823 876 826
rect 1274 816 1277 825
rect 1378 816 1381 825
rect 1450 823 1461 826
rect 1450 816 1453 823
rect 1922 816 1925 825
rect 2490 823 2500 826
rect 2530 823 2548 826
rect 340 813 357 816
rect 372 813 381 816
rect 420 813 437 816
rect 556 813 565 816
rect 596 813 605 816
rect 652 813 661 816
rect 706 813 716 816
rect 892 813 908 816
rect 914 813 924 816
rect 954 813 980 816
rect 1058 813 1068 816
rect 1074 813 1084 816
rect 1114 813 1140 816
rect 1204 813 1228 816
rect 1242 813 1260 816
rect 1274 813 1285 816
rect 1300 813 1324 816
rect 1346 813 1356 816
rect 1370 813 1381 816
rect 164 803 172 806
rect 316 803 333 806
rect 428 803 452 806
rect 474 803 492 806
rect 658 805 661 813
rect 684 803 701 806
rect 914 805 917 813
rect 1058 806 1061 813
rect 1044 803 1061 806
rect 1074 805 1077 813
rect 1178 803 1196 806
rect 1018 793 1028 796
rect 1282 795 1285 813
rect 1292 803 1309 806
rect 1332 803 1348 806
rect 1370 805 1373 813
rect 1410 805 1413 816
rect 1444 813 1453 816
rect 1458 813 1468 816
rect 1474 805 1477 816
rect 1482 813 1492 816
rect 1554 813 1580 816
rect 1652 813 1661 816
rect 1708 813 1717 816
rect 1722 805 1725 816
rect 1762 813 1772 816
rect 1762 806 1765 813
rect 1756 803 1765 806
rect 1778 805 1781 816
rect 1898 813 1908 816
rect 1922 813 1940 816
rect 2172 813 2212 816
rect 2356 813 2373 816
rect 2516 813 2549 816
rect 2698 813 2725 816
rect 1924 803 1933 806
rect 1948 803 1973 806
rect 2098 803 2108 806
rect 2330 803 2348 806
rect 2362 803 2372 806
rect 2490 803 2500 806
rect 2684 803 2701 806
rect 2722 805 2725 813
rect 2746 813 2781 816
rect 2852 813 2861 816
rect 2866 813 2876 816
rect 2890 813 2901 816
rect 2746 805 2749 813
rect 2812 803 2837 806
rect 2890 805 2893 813
rect 2946 803 2949 814
rect 2978 813 2996 816
rect 2970 803 2988 806
rect 2754 793 2804 796
rect 38 767 3053 773
rect 3871 767 3889 1061
rect 4601 864 4650 911
rect 3871 761 3900 767
rect 330 743 340 746
rect 1164 743 1173 746
rect 170 726 173 735
rect 324 733 341 736
rect 348 733 365 736
rect 482 733 500 736
rect 530 733 540 736
rect 554 733 564 736
rect 692 733 725 736
rect 900 733 909 736
rect 1026 733 1036 736
rect 1140 733 1156 736
rect 1162 733 1180 736
rect 108 723 133 726
rect 164 723 173 726
rect 308 723 317 726
rect 332 723 341 726
rect 362 725 365 733
rect 1026 726 1029 733
rect 1186 726 1189 745
rect 1282 743 1292 746
rect 1218 733 1236 736
rect 1276 733 1293 736
rect 460 723 469 726
rect 508 723 517 726
rect 524 723 541 726
rect 548 723 572 726
rect 604 723 621 726
rect 658 723 676 726
rect 756 723 765 726
rect 1020 723 1029 726
rect 1090 723 1108 726
rect 1186 723 1213 726
rect 1244 723 1253 726
rect 1308 723 1316 726
rect 1460 723 1485 726
rect 1522 725 1525 736
rect 1540 733 1564 736
rect 1698 726 1701 735
rect 1946 733 1988 736
rect 2012 733 2037 736
rect 2154 726 2157 735
rect 2282 733 2300 736
rect 2348 733 2365 736
rect 2370 733 2380 736
rect 2498 726 2501 735
rect 2642 726 2645 735
rect 2714 733 2724 736
rect 2802 733 2820 736
rect 2842 733 2868 736
rect 2892 733 2909 736
rect 2948 733 2980 736
rect 1580 723 1597 726
rect 1692 723 1701 726
rect 1724 723 1733 726
rect 1780 723 1805 726
rect 1874 723 1892 726
rect 1906 723 1924 726
rect 1978 723 1996 726
rect 2092 723 2117 726
rect 2148 723 2157 726
rect 2164 723 2173 726
rect 2218 723 2244 726
rect 2282 723 2308 726
rect 2322 723 2340 726
rect 2436 723 2461 726
rect 2492 723 2501 726
rect 2636 723 2645 726
rect 2658 723 2684 726
rect 2714 723 2732 726
rect 2762 723 2772 726
rect 2842 725 2845 733
rect 2850 723 2876 726
rect 2898 723 2924 726
rect 588 713 597 716
rect 652 713 661 716
rect 692 713 701 716
rect 1116 713 1124 716
rect 1906 715 1909 723
rect 2322 715 2325 723
rect 3871 718 3889 761
rect 410 703 436 706
rect 618 703 644 706
rect 14 667 3077 673
rect 418 633 444 636
rect 2418 626 2421 636
rect 3900 626 3908 631
rect 394 623 404 626
rect 428 623 437 626
rect 636 623 645 626
rect 890 623 908 626
rect 2266 616 2269 625
rect 2412 623 2421 626
rect 2506 623 2548 626
rect 2634 623 2676 626
rect 3892 621 3908 626
rect 3884 616 3908 621
rect 116 613 141 616
rect 172 613 181 616
rect 252 613 269 616
rect 298 613 324 616
rect 354 613 364 616
rect 370 613 405 616
rect 412 613 421 616
rect 468 613 477 616
rect 178 605 181 613
rect 234 603 244 606
rect 292 603 317 606
rect 354 596 357 613
rect 370 605 373 613
rect 522 606 525 614
rect 564 613 573 616
rect 580 613 620 616
rect 652 613 669 616
rect 690 613 701 616
rect 740 613 773 616
rect 924 613 933 616
rect 1042 613 1060 616
rect 1090 613 1108 616
rect 1170 613 1196 616
rect 1252 613 1268 616
rect 1332 613 1349 616
rect 1394 613 1404 616
rect 1484 613 1500 616
rect 1540 613 1548 616
rect 1578 613 1588 616
rect 1700 613 1709 616
rect 1772 613 1781 616
rect 1884 613 1901 616
rect 1938 613 1956 616
rect 2066 613 2076 616
rect 2116 613 2125 616
rect 2220 613 2229 616
rect 2236 613 2252 616
rect 2266 613 2284 616
rect 2404 613 2421 616
rect 2428 613 2445 616
rect 2452 613 2485 616
rect 2570 613 2661 616
rect 2698 613 2716 616
rect 2730 613 2740 616
rect 2770 613 2796 616
rect 2938 613 2996 616
rect 396 603 405 606
rect 492 603 508 606
rect 522 603 556 606
rect 594 603 612 606
rect 658 603 668 606
rect 690 605 693 613
rect 748 603 773 606
rect 884 603 901 606
rect 1090 603 1100 606
rect 1338 603 1348 606
rect 1452 603 1461 606
rect 1738 603 1748 606
rect 1780 603 1789 606
rect 1898 605 1901 613
rect 1940 603 1949 606
rect 2226 605 2229 613
rect 2268 603 2277 606
rect 2410 603 2420 606
rect 2434 603 2444 606
rect 2500 603 2541 606
rect 2570 605 2573 613
rect 2628 603 2661 606
rect 2698 605 2701 613
rect 2730 606 2733 613
rect 3876 610 3908 616
rect 2724 603 2733 606
rect 2842 603 2860 606
rect 2940 603 2988 606
rect 194 593 220 596
rect 348 593 357 596
rect 38 567 3053 573
rect 3128 565 3908 610
rect 300 543 308 546
rect 122 533 132 536
rect 226 533 236 536
rect 292 533 309 536
rect 330 533 372 536
rect 386 533 396 536
rect 444 533 468 536
rect 482 533 500 536
rect 578 533 596 536
rect 1156 533 1164 536
rect 1364 533 1373 536
rect 1410 533 1428 536
rect 226 526 229 533
rect 162 523 229 526
rect 274 523 284 526
rect 380 523 397 526
rect 404 523 421 526
rect 476 523 493 526
rect 572 523 597 526
rect 412 513 428 516
rect 532 513 541 516
rect 556 513 565 516
rect 580 513 589 516
rect 620 513 629 516
rect 658 513 668 516
rect 674 506 677 525
rect 740 523 749 526
rect 780 523 812 526
rect 818 523 828 526
rect 1034 523 1044 526
rect 1124 523 1148 526
rect 1162 523 1172 526
rect 1260 523 1285 526
rect 1346 523 1356 526
rect 1410 516 1413 533
rect 1418 523 1436 526
rect 1450 523 1453 534
rect 1532 533 1549 536
rect 1612 533 1637 536
rect 1738 533 1748 536
rect 1828 533 1837 536
rect 2234 526 2237 534
rect 2394 533 2404 536
rect 2674 533 2692 536
rect 2708 533 2756 536
rect 2786 533 2796 536
rect 2674 526 2677 533
rect 1474 523 1508 526
rect 1562 523 1572 526
rect 1578 523 1596 526
rect 1756 523 1780 526
rect 1860 523 1868 526
rect 2068 523 2092 526
rect 2124 523 2133 526
rect 2228 523 2237 526
rect 2244 523 2260 526
rect 2388 523 2405 526
rect 2412 523 2421 526
rect 2660 523 2677 526
rect 2716 523 2764 526
rect 2786 523 2804 526
rect 2842 525 2845 536
rect 2852 533 2877 536
rect 2906 526 2909 534
rect 2906 523 2917 526
rect 2938 523 2948 526
rect 2786 516 2789 523
rect 692 513 701 516
rect 722 513 732 516
rect 1082 513 1108 516
rect 1370 513 1380 516
rect 1404 513 1413 516
rect 1476 513 1493 516
rect 1612 513 1621 516
rect 2722 513 2741 516
rect 2780 513 2789 516
rect 2914 515 2917 523
rect 530 503 548 506
rect 666 503 677 506
rect 1388 503 1397 506
rect 14 467 3077 473
rect -144 391 58 436
rect 1492 433 1517 436
rect 404 423 413 426
rect 484 423 492 426
rect 658 423 668 426
rect 1452 423 1461 426
rect 148 413 157 416
rect 194 413 228 416
rect 236 413 277 416
rect 372 413 381 416
rect 396 413 429 416
rect 436 413 453 416
rect 476 413 493 416
rect 500 413 509 416
rect 652 413 669 416
rect 722 413 732 416
rect 780 413 789 416
rect 1212 413 1220 416
rect 1324 413 1333 416
rect 196 403 213 406
rect 244 403 261 406
rect 274 395 277 413
rect 308 403 325 406
rect 332 403 364 406
rect 402 403 428 406
rect 450 403 453 413
rect 610 403 644 406
rect 1386 403 1389 414
rect 1402 413 1412 416
rect 316 393 324 396
rect 1402 395 1405 413
rect 1434 403 1437 414
rect 1468 413 1477 416
rect 1514 405 1517 433
rect 1562 416 1565 425
rect 2242 416 2245 425
rect 2292 423 2300 426
rect 2562 423 2580 426
rect 2922 416 2925 425
rect 2956 423 2965 426
rect 1524 413 1541 416
rect 1562 413 1573 416
rect 1620 413 1637 416
rect 1652 413 1677 416
rect 1812 413 1852 416
rect 1972 413 1997 416
rect 2028 413 2037 416
rect 2204 413 2213 416
rect 2218 413 2228 416
rect 2242 413 2260 416
rect 2436 413 2461 416
rect 2602 413 2676 416
rect 2812 413 2837 416
rect 2882 413 2892 416
rect 2898 413 2916 416
rect 2922 413 2940 416
rect 1570 405 1573 413
rect 1596 403 1605 406
rect 1626 403 1636 406
rect 1786 403 1804 406
rect 1818 403 1844 406
rect 2034 403 2044 406
rect 2266 403 2276 406
rect 2418 403 2428 406
rect 2602 405 2605 413
rect 2700 403 2709 406
rect 2754 403 2804 406
rect 2818 403 2836 406
rect 2860 403 2885 406
rect 2898 405 2901 413
rect 2922 403 2932 406
rect 38 367 3053 373
rect 468 333 485 336
rect 674 333 684 336
rect 794 333 812 336
rect 108 323 133 326
rect 260 323 276 326
rect 492 323 501 326
rect 580 323 605 326
rect 652 323 660 326
rect 972 323 1004 326
rect 1010 323 1020 326
rect 1052 323 1068 326
rect 1074 323 1084 326
rect 1114 323 1140 326
rect 1234 323 1237 334
rect 1338 326 1341 334
rect 1564 333 1580 336
rect 1332 323 1341 326
rect 1354 323 1372 326
rect 1500 323 1509 326
rect 1524 323 1541 326
rect 1546 323 1556 326
rect 1602 323 1605 334
rect 1884 333 1900 336
rect 2074 326 2077 334
rect 2202 333 2252 336
rect 2276 333 2285 336
rect 2308 333 2317 336
rect 2434 333 2444 336
rect 2506 326 2509 334
rect 2964 333 2973 336
rect 1612 323 1621 326
rect 1876 323 1901 326
rect 2012 323 2037 326
rect 2068 323 2077 326
rect 2132 323 2157 326
rect 2188 323 2197 326
rect 2202 323 2260 326
rect 2282 323 2300 326
rect 2428 323 2445 326
rect 2452 323 2477 326
rect 2506 323 2533 326
rect 2572 323 2581 326
rect 2690 323 2708 326
rect 2714 323 2732 326
rect 2874 323 2884 326
rect 498 316 501 323
rect 2282 316 2285 323
rect 498 313 517 316
rect 532 313 541 316
rect 594 313 612 316
rect 788 313 805 316
rect 1420 313 1428 316
rect 1538 313 1548 316
rect 1634 313 1644 316
rect 2276 313 2285 316
rect 2474 316 2477 323
rect 2474 313 2484 316
rect 2650 313 2668 316
rect 498 303 524 306
rect 586 303 628 306
rect 1466 303 1476 306
rect 2906 303 2924 306
rect 14 267 3077 273
rect 522 233 540 236
rect 1594 233 1604 236
rect 524 223 533 226
rect 548 223 557 226
rect 684 223 693 226
rect 754 216 757 225
rect 924 223 957 226
rect 1428 223 1436 226
rect 1546 223 1556 226
rect 1634 223 1645 226
rect 1634 216 1637 223
rect 2146 216 2149 225
rect 2226 216 2229 225
rect 2650 223 2676 226
rect 3128 225 3173 565
rect 2938 216 2941 225
rect 108 213 133 216
rect 196 213 205 216
rect 242 213 252 216
rect 354 213 413 216
rect 436 213 453 216
rect 580 213 589 216
rect 626 213 637 216
rect 644 213 661 216
rect 668 213 677 216
rect 276 203 293 206
rect 314 203 324 206
rect 354 205 357 213
rect 372 203 389 206
rect 282 193 292 196
rect 402 193 412 196
rect 450 195 453 213
rect 474 203 500 206
rect 626 205 629 213
rect 634 205 637 213
rect 650 203 660 206
rect 690 203 693 214
rect 730 213 741 216
rect 754 214 764 216
rect 754 213 765 214
rect 852 213 877 216
rect 988 213 997 216
rect 738 205 741 213
rect 762 203 765 213
rect 866 203 876 206
rect 946 203 964 206
rect 1106 205 1109 216
rect 1242 205 1245 216
rect 1340 213 1349 216
rect 1356 213 1380 216
rect 1346 205 1349 213
rect 1362 203 1372 206
rect 1410 203 1413 214
rect 1476 213 1493 216
rect 1620 213 1637 216
rect 1820 213 1845 216
rect 1876 213 1885 216
rect 1562 203 1572 206
rect 1628 203 1637 206
rect 1898 205 1901 216
rect 1980 213 1997 216
rect 2092 213 2101 216
rect 2108 213 2132 216
rect 2146 213 2164 216
rect 2170 213 2212 216
rect 2226 213 2244 216
rect 2250 213 2300 216
rect 2338 213 2356 216
rect 2460 213 2469 216
rect 2484 213 2501 216
rect 2698 213 2724 216
rect 2844 213 2853 216
rect 2866 213 2876 216
rect 2908 213 2917 216
rect 2938 213 2948 216
rect 2098 205 2101 213
rect 2466 206 2469 213
rect 2178 203 2204 206
rect 2252 203 2277 206
rect 2316 203 2325 206
rect 2340 203 2349 206
rect 2466 203 2476 206
rect 2490 203 2500 206
rect 2700 203 2709 206
rect 2850 205 2853 213
rect 2884 203 2893 206
rect 2914 205 2917 213
rect 2956 203 2973 206
rect 3033 180 3173 225
rect 38 167 3053 173
rect 252 143 260 146
rect 442 143 452 146
rect 186 126 189 134
rect 244 133 261 136
rect 268 133 293 136
rect 436 133 453 136
rect 460 133 493 136
rect 498 133 508 136
rect 570 133 596 136
rect 618 126 621 134
rect 634 133 652 136
rect 682 126 685 145
rect 1378 143 1388 146
rect 692 133 701 136
rect 706 133 724 136
rect 842 133 860 136
rect 116 123 141 126
rect 172 123 189 126
rect 196 123 236 126
rect 332 123 341 126
rect 474 123 500 126
rect 538 123 556 126
rect 562 123 621 126
rect 628 123 645 126
rect 676 123 685 126
rect 732 123 757 126
rect 778 123 788 126
rect 882 125 885 136
rect 906 133 924 136
rect 972 133 989 136
rect 1210 126 1213 134
rect 1372 133 1381 136
rect 948 123 964 126
rect 1132 123 1141 126
rect 1188 123 1213 126
rect 1324 123 1333 126
rect 1380 123 1389 126
rect 1418 125 1421 136
rect 1458 133 1468 136
rect 1482 133 1516 136
rect 1970 126 1973 134
rect 2290 133 2300 136
rect 2324 133 2333 136
rect 2434 133 2444 136
rect 2458 133 2468 136
rect 2434 126 2437 133
rect 2618 126 2621 134
rect 2700 133 2709 136
rect 2938 133 2948 136
rect 1442 123 1452 126
rect 1466 123 1476 126
rect 1524 123 1572 126
rect 1812 123 1837 126
rect 1908 123 1933 126
rect 1964 123 1973 126
rect 1980 123 2069 126
rect 2108 123 2133 126
rect 2164 123 2173 126
rect 2220 123 2229 126
rect 2282 123 2308 126
rect 2428 123 2437 126
rect 2452 123 2469 126
rect 2612 123 2621 126
rect 2804 123 2813 126
rect 2820 123 2837 126
rect 2922 123 2932 126
rect 2938 123 2956 126
rect 564 113 573 116
rect 740 113 764 116
rect 876 113 885 116
rect 900 113 917 116
rect 1436 113 1445 116
rect 1532 113 1557 116
rect 2634 113 2676 116
rect 2892 113 2901 116
rect 2916 113 2925 116
rect 2938 115 2941 123
rect 874 103 892 106
rect 1410 103 1428 106
rect 2882 103 2908 106
rect 14 67 3077 73
rect 38 37 3053 57
rect 14 13 3077 33
rect 441 -30 497 13
rect -851 -48 497 -30
rect -851 -133 -839 -48
rect -862 -139 -839 -133
rect -1608 -338 -1571 -291
rect -823 -433 -805 -70
rect -862 -439 -805 -433
rect -1605 -633 -1566 -585
rect -823 -701 -805 -439
rect -823 -719 350 -701
rect -823 -727 -817 -719
rect -865 -733 -817 -727
rect -852 -737 -817 -733
rect -852 -743 -846 -737
rect -558 -743 -552 -719
rect -258 -743 -251 -719
rect 42 -725 48 -719
rect 441 -726 497 -48
rect 2109 -701 2145 -692
rect 560 -707 2145 -701
rect 560 -716 2136 -707
rect 560 -719 2127 -716
rect 2241 -717 2297 13
rect 3847 -692 3862 565
rect 3876 560 3908 565
rect 3884 555 3908 560
rect 4603 558 4644 617
rect 3892 550 3908 555
rect 3900 545 3908 550
rect 2441 -707 3862 -692
rect 3871 167 3889 457
rect 4611 260 4646 311
rect 3871 161 3900 167
rect 3871 -133 3889 161
rect 4612 -35 4645 10
rect 3871 -139 3900 -133
rect 3871 -433 3889 -139
rect 4609 -341 4645 -283
rect 3871 -439 3900 -433
rect 2241 -719 2751 -717
rect 3871 -719 3889 -439
rect 4605 -641 4649 -588
rect 642 -725 648 -719
rect 942 -725 948 -719
rect 1242 -725 1248 -719
rect 1542 -725 1548 -719
rect 1842 -725 1848 -719
rect 2241 -721 3889 -719
rect 2241 -723 3890 -721
rect 2241 -724 3891 -723
rect 2241 -725 3892 -724
rect 2241 -726 3893 -725
rect 436 -734 502 -726
rect 2236 -734 2302 -726
rect 2742 -727 3894 -726
rect 2742 -728 3895 -727
rect 2742 -729 3896 -728
rect 2742 -730 3883 -729
rect 3886 -730 3896 -729
rect 2742 -731 3882 -730
rect 3887 -731 3897 -730
rect 2742 -733 3881 -731
rect 3888 -732 3898 -731
rect 3889 -733 3899 -732
rect 2742 -734 3880 -733
rect 3890 -734 3900 -733
rect 431 -742 507 -734
rect 2231 -742 2307 -734
rect 426 -750 512 -742
rect 2226 -750 2312 -742
rect 2742 -743 2748 -734
rect 3042 -743 3048 -734
rect 3342 -743 3348 -734
rect 3642 -743 3648 -734
rect 3891 -736 3900 -734
rect 3892 -738 3900 -736
rect 3894 -739 3900 -738
rect -758 -1486 -705 -1448
rect -452 -1485 -411 -1454
rect -147 -1485 -114 -1455
rect 435 -1487 501 -1447
rect 2231 -1495 2310 -1451
rect 2539 -1496 2599 -1449
rect 2842 -1493 2900 -1454
rect 3142 -1496 3202 -1453
rect 3442 -1497 3498 -1448
rect 3740 -1489 3798 -1450
<< metal2 >>
rect -858 4013 -852 4019
rect -835 3810 -830 4019
rect -558 4013 -552 4019
rect -535 3836 -530 4019
rect -258 4013 -252 4019
rect -235 3855 -230 4019
rect 42 4013 48 4019
rect -235 3850 32 3855
rect -535 3831 12 3836
rect -835 3805 -15 3810
rect -862 3784 -38 3789
rect -862 3761 -856 3767
rect -862 3697 -56 3702
rect -862 3461 -823 3467
rect -862 3397 -74 3402
rect -79 3239 -74 3397
rect -61 3271 -56 3697
rect -43 3298 -38 3784
rect -20 3324 -15 3805
rect 7 3352 12 3831
rect 27 3372 32 3850
rect 65 3400 70 4019
rect 342 3980 348 4019
rect 578 3426 583 4019
rect 642 3980 648 4019
rect 878 3455 883 4019
rect 1242 3980 1248 4019
rect 942 3962 1196 3980
rect 1478 3484 1483 4019
rect 1542 4013 1548 4019
rect 1565 3505 1570 4019
rect 1842 4013 1848 4019
rect 1865 3536 1870 4019
rect 2142 4013 2148 4019
rect 2165 3952 2170 4019
rect 2442 4013 2448 4019
rect 2015 3947 2170 3952
rect 1865 3531 1926 3536
rect 1565 3500 1854 3505
rect 1478 3479 1599 3484
rect 878 3450 1581 3455
rect 578 3421 1534 3426
rect 65 3395 1520 3400
rect 27 3367 1504 3372
rect 7 3347 1477 3352
rect -20 3319 1462 3324
rect -43 3293 1382 3298
rect -61 3266 1303 3271
rect -79 3234 1238 3239
rect -79 3206 1166 3211
rect -862 3161 -823 3167
rect -79 3102 -74 3206
rect -862 3097 -74 3102
rect -66 3186 862 3191
rect -862 2861 -823 2867
rect -851 2552 -839 2822
rect -66 2590 -61 3186
rect -139 2585 -61 2590
rect -53 3153 838 3158
rect -862 2509 -856 2515
rect -139 2492 -134 2585
rect -53 2564 -48 3153
rect -862 2487 -134 2492
rect -126 2559 -48 2564
rect -40 3122 750 3127
rect -126 1989 -121 2559
rect -40 2531 -35 3122
rect -862 1984 -121 1989
rect -113 2526 -35 2531
rect -27 3092 607 3097
rect -862 1961 -856 1967
rect -113 1689 -108 2526
rect -27 2489 -22 3092
rect -862 1684 -108 1689
rect -100 2484 -22 2489
rect -13 3065 478 3070
rect -862 1661 -856 1667
rect -100 1602 -95 2484
rect -13 2453 -8 3065
rect -862 1597 -95 1602
rect -87 2448 -8 2453
rect 2 3040 326 3045
rect 473 3040 478 3065
rect 602 3040 607 3092
rect 745 3040 750 3122
rect 833 3040 838 3153
rect 857 3040 862 3186
rect 1161 3040 1166 3206
rect 1233 3040 1238 3234
rect 1298 3045 1303 3266
rect 1297 3040 1303 3045
rect 1377 3040 1382 3293
rect 1457 3040 1462 3319
rect 1472 3051 1477 3347
rect 1499 3051 1504 3367
rect 1472 3046 1478 3051
rect 1473 3040 1478 3046
rect 1497 3046 1504 3051
rect 1515 3049 1520 3395
rect 1497 3040 1502 3046
rect 1513 3044 1520 3049
rect 1513 3040 1518 3044
rect 1529 3040 1534 3421
rect 1576 3051 1581 3450
rect 1594 3061 1599 3479
rect 1593 3056 1599 3061
rect 1576 3046 1582 3051
rect 1577 3040 1582 3046
rect 1593 3040 1598 3056
rect 1849 3040 1854 3500
rect 1921 3040 1926 3531
rect 2015 3040 2020 3947
rect 2465 3213 2470 4019
rect 2742 4013 2748 4019
rect 2102 3208 2470 3213
rect 2102 3059 2107 3208
rect 2765 3194 2770 4019
rect 3342 4013 3348 4019
rect 3040 3962 3289 3980
rect 2097 3054 2107 3059
rect 2146 3189 2770 3194
rect 2097 3040 2102 3054
rect 2146 3053 2151 3189
rect 3365 3178 3370 4019
rect 3642 4013 3648 4019
rect 2263 3173 3370 3178
rect 2263 3105 2268 3173
rect 3665 3160 3670 4019
rect 2145 3048 2151 3053
rect 2262 3100 2268 3105
rect 2279 3155 3670 3160
rect 3684 3784 3900 3789
rect 2262 3050 2267 3100
rect 2145 3040 2150 3048
rect 2262 3045 2270 3050
rect 2265 3040 2270 3045
rect 2279 3047 2284 3155
rect 3684 3146 3689 3784
rect 3894 3761 3900 3767
rect 2417 3141 3689 3146
rect 3706 3484 3900 3489
rect 2417 3081 2422 3141
rect 3706 3132 3711 3484
rect 3894 3461 3900 3467
rect 2416 3076 2422 3081
rect 2441 3127 3711 3132
rect 3729 3184 3900 3189
rect 2279 3042 2286 3047
rect 2281 3040 2286 3042
rect 2416 3040 2421 3076
rect 2441 3040 2446 3127
rect 3729 3112 3734 3184
rect 3894 3161 3900 3167
rect 2641 3107 3734 3112
rect 2641 3040 2646 3107
rect 2752 3087 3854 3092
rect 2752 3050 2757 3087
rect 2816 3059 3822 3064
rect 2752 3045 2758 3050
rect 2753 3040 2758 3045
rect 2816 3045 2821 3059
rect 2816 3040 2822 3045
rect -862 1361 -823 1367
rect -87 1302 -82 2448
rect 2 2404 7 3040
rect -862 1297 -82 1302
rect -74 2399 7 2404
rect -862 1061 -823 1067
rect -851 755 -839 1031
rect -74 479 -69 2399
rect -862 474 -69 479
rect -62 2362 0 2367
rect -862 184 -821 189
rect -62 184 -57 2362
rect -826 179 -57 184
rect -50 2292 0 2297
rect -862 161 -856 167
rect -50 102 -45 2292
rect -23 2012 -1 2017
rect -23 1959 -18 2012
rect -135 97 -45 102
rect -38 1954 -18 1959
rect -823 -88 -805 15
rect -862 -116 -830 -111
rect -835 -117 -830 -116
rect -135 -117 -130 97
rect -38 82 -33 1954
rect -6 1942 -1 1997
rect -835 -122 -130 -117
rect -112 77 -33 82
rect -26 1937 -1 1942
rect -862 -139 -856 -133
rect -112 -198 -107 77
rect -26 58 -21 1937
rect -862 -203 -107 -198
rect -83 53 -21 58
rect -15 1922 0 1927
rect -862 -439 -856 -433
rect -83 -498 -78 53
rect -15 27 -10 1922
rect -862 -503 -78 -498
rect -61 22 -10 27
rect -61 -654 -56 22
rect -5 8 0 1907
rect 14 13 34 3027
rect 38 37 58 3003
rect 322 2966 325 3040
rect 314 2963 325 2966
rect 82 2523 85 2926
rect 122 2923 125 2936
rect 314 2933 317 2963
rect 170 2843 173 2926
rect 186 2923 205 2926
rect 218 2923 261 2926
rect 114 2503 117 2836
rect 138 2833 157 2836
rect 122 2723 125 2826
rect 130 2813 133 2826
rect 146 2813 149 2826
rect 154 2823 157 2833
rect 162 2756 165 2826
rect 170 2806 173 2836
rect 178 2823 181 2836
rect 186 2806 189 2923
rect 234 2896 237 2916
rect 242 2913 253 2916
rect 258 2913 261 2923
rect 242 2903 261 2906
rect 234 2893 245 2896
rect 170 2803 189 2806
rect 194 2803 197 2816
rect 202 2803 205 2816
rect 210 2766 213 2846
rect 234 2793 237 2816
rect 206 2763 213 2766
rect 154 2753 165 2756
rect 130 2733 149 2736
rect 130 2703 133 2733
rect 154 2726 157 2753
rect 170 2733 173 2746
rect 186 2743 189 2756
rect 146 2723 157 2726
rect 138 2683 141 2716
rect 154 2713 157 2723
rect 170 2696 173 2726
rect 186 2723 189 2736
rect 194 2723 197 2736
rect 206 2716 209 2763
rect 242 2733 245 2893
rect 258 2833 261 2903
rect 250 2823 261 2826
rect 266 2823 269 2926
rect 314 2913 317 2926
rect 162 2693 173 2696
rect 162 2636 165 2693
rect 162 2633 173 2636
rect 130 2593 133 2616
rect 170 2613 173 2633
rect 178 2613 181 2716
rect 206 2713 213 2716
rect 210 2693 213 2713
rect 242 2706 245 2726
rect 234 2703 245 2706
rect 234 2636 237 2703
rect 234 2633 245 2636
rect 130 2523 133 2546
rect 186 2533 189 2606
rect 194 2533 197 2616
rect 210 2613 213 2626
rect 202 2593 205 2606
rect 202 2533 205 2546
rect 66 2343 69 2406
rect 130 2403 133 2416
rect 66 2213 69 2336
rect 90 2333 117 2336
rect 122 2333 133 2336
rect 114 2273 117 2326
rect 122 2213 125 2333
rect 130 2323 149 2326
rect 130 2303 133 2316
rect 154 2193 157 2526
rect 186 2503 189 2526
rect 194 2513 197 2526
rect 210 2503 213 2526
rect 218 2516 221 2606
rect 226 2523 229 2606
rect 234 2596 237 2616
rect 242 2603 245 2633
rect 250 2613 253 2823
rect 266 2803 269 2816
rect 274 2743 277 2836
rect 290 2793 293 2836
rect 274 2663 277 2736
rect 290 2703 293 2756
rect 274 2613 277 2626
rect 234 2593 261 2596
rect 266 2593 269 2606
rect 282 2603 285 2696
rect 298 2623 301 2806
rect 314 2803 317 2826
rect 322 2803 325 2956
rect 330 2846 333 2916
rect 338 2883 341 2936
rect 354 2903 357 2926
rect 330 2843 341 2846
rect 338 2813 341 2843
rect 322 2743 325 2796
rect 338 2736 341 2806
rect 346 2753 349 2826
rect 362 2816 365 2936
rect 354 2813 365 2816
rect 370 2813 373 2826
rect 306 2703 309 2726
rect 330 2723 333 2736
rect 338 2733 349 2736
rect 314 2666 317 2716
rect 338 2703 341 2726
rect 314 2663 325 2666
rect 234 2516 237 2526
rect 242 2523 245 2536
rect 218 2513 237 2516
rect 234 2436 237 2513
rect 194 2416 197 2426
rect 202 2423 213 2426
rect 170 2376 173 2406
rect 162 2373 173 2376
rect 162 2316 165 2373
rect 170 2333 173 2356
rect 178 2323 181 2416
rect 194 2413 205 2416
rect 186 2403 197 2406
rect 162 2313 189 2316
rect 194 2306 197 2396
rect 202 2316 205 2413
rect 210 2393 213 2423
rect 218 2413 221 2436
rect 234 2433 245 2436
rect 250 2433 253 2526
rect 258 2436 261 2593
rect 298 2583 301 2606
rect 258 2433 269 2436
rect 242 2426 245 2433
rect 234 2373 237 2426
rect 242 2423 253 2426
rect 242 2393 245 2406
rect 210 2323 221 2326
rect 202 2313 213 2316
rect 218 2313 221 2323
rect 234 2313 237 2326
rect 194 2303 205 2306
rect 242 2303 245 2346
rect 250 2313 253 2423
rect 258 2413 261 2426
rect 266 2396 269 2433
rect 258 2393 269 2396
rect 258 2346 261 2366
rect 266 2356 269 2393
rect 274 2426 277 2446
rect 282 2433 285 2526
rect 274 2423 285 2426
rect 274 2363 277 2423
rect 282 2413 285 2423
rect 290 2413 293 2426
rect 306 2406 309 2616
rect 314 2603 317 2616
rect 322 2613 325 2663
rect 346 2636 349 2733
rect 354 2643 357 2813
rect 362 2793 365 2806
rect 386 2803 389 2886
rect 394 2823 397 2926
rect 402 2913 413 2916
rect 394 2796 397 2816
rect 402 2803 405 2836
rect 410 2813 413 2826
rect 410 2796 413 2806
rect 394 2793 413 2796
rect 418 2786 421 2936
rect 458 2916 461 2936
rect 474 2933 477 3040
rect 602 2986 605 3040
rect 602 2983 621 2986
rect 522 2926 525 2966
rect 530 2933 533 2946
rect 538 2933 541 2956
rect 602 2936 605 2976
rect 570 2933 581 2936
rect 586 2933 605 2936
rect 610 2933 613 2946
rect 514 2923 525 2926
rect 450 2913 461 2916
rect 450 2846 453 2913
rect 450 2843 461 2846
rect 458 2826 461 2843
rect 426 2806 429 2816
rect 434 2813 445 2816
rect 426 2803 437 2806
rect 434 2793 437 2803
rect 410 2783 421 2786
rect 362 2733 365 2756
rect 362 2703 365 2726
rect 370 2723 373 2736
rect 346 2633 357 2636
rect 330 2623 349 2626
rect 330 2603 333 2623
rect 338 2603 341 2616
rect 346 2613 349 2623
rect 346 2593 349 2606
rect 354 2603 357 2633
rect 370 2606 373 2616
rect 362 2603 373 2606
rect 362 2523 365 2603
rect 378 2593 381 2746
rect 386 2733 389 2756
rect 402 2733 405 2756
rect 386 2693 389 2726
rect 402 2703 405 2726
rect 402 2603 405 2626
rect 410 2606 413 2783
rect 442 2746 445 2813
rect 450 2753 453 2826
rect 458 2823 469 2826
rect 474 2823 477 2916
rect 506 2903 509 2916
rect 458 2803 461 2816
rect 466 2746 469 2823
rect 418 2743 429 2746
rect 434 2743 445 2746
rect 462 2743 469 2746
rect 426 2706 429 2726
rect 422 2703 429 2706
rect 422 2626 425 2703
rect 422 2623 429 2626
rect 410 2603 421 2606
rect 426 2603 429 2623
rect 434 2613 437 2743
rect 442 2713 445 2736
rect 442 2673 445 2706
rect 450 2703 453 2726
rect 462 2696 465 2743
rect 474 2723 477 2736
rect 482 2723 485 2816
rect 498 2803 501 2816
rect 506 2786 509 2826
rect 522 2813 525 2826
rect 538 2823 541 2926
rect 562 2913 565 2926
rect 570 2923 581 2926
rect 594 2913 597 2926
rect 618 2916 621 2983
rect 610 2913 621 2916
rect 502 2783 509 2786
rect 490 2703 493 2716
rect 502 2706 505 2783
rect 502 2703 509 2706
rect 450 2693 465 2696
rect 442 2613 445 2626
rect 450 2603 453 2693
rect 410 2583 413 2596
rect 418 2593 421 2603
rect 466 2583 469 2596
rect 386 2533 389 2546
rect 314 2413 317 2426
rect 322 2413 325 2436
rect 362 2426 365 2516
rect 402 2513 405 2526
rect 338 2413 341 2426
rect 362 2423 373 2426
rect 354 2413 365 2416
rect 282 2393 285 2406
rect 266 2353 277 2356
rect 258 2343 269 2346
rect 258 2313 261 2326
rect 266 2303 269 2343
rect 274 2333 277 2353
rect 290 2333 293 2406
rect 306 2403 317 2406
rect 322 2333 325 2346
rect 330 2333 333 2406
rect 338 2393 341 2406
rect 346 2393 349 2406
rect 370 2403 373 2423
rect 282 2313 285 2326
rect 186 2193 189 2206
rect 234 2193 237 2216
rect 274 2213 277 2256
rect 290 2223 293 2326
rect 290 2213 309 2216
rect 314 2213 317 2326
rect 322 2313 325 2326
rect 330 2223 333 2266
rect 338 2213 341 2326
rect 354 2303 357 2316
rect 346 2223 349 2236
rect 354 2206 357 2226
rect 362 2213 365 2346
rect 370 2263 373 2316
rect 378 2303 381 2436
rect 418 2416 421 2526
rect 474 2523 477 2616
rect 490 2603 493 2696
rect 506 2683 509 2703
rect 514 2686 517 2756
rect 522 2713 525 2806
rect 530 2793 533 2816
rect 538 2803 541 2816
rect 554 2813 557 2826
rect 562 2813 565 2906
rect 610 2836 613 2913
rect 610 2833 621 2836
rect 530 2716 533 2736
rect 538 2733 541 2776
rect 562 2756 565 2806
rect 570 2773 573 2826
rect 578 2813 589 2816
rect 562 2753 573 2756
rect 554 2723 557 2736
rect 530 2713 549 2716
rect 562 2713 565 2736
rect 570 2733 573 2753
rect 578 2723 581 2736
rect 586 2723 589 2806
rect 514 2683 525 2686
rect 514 2616 517 2626
rect 506 2613 517 2616
rect 506 2533 509 2546
rect 522 2533 525 2683
rect 530 2596 533 2636
rect 546 2633 549 2713
rect 538 2616 541 2626
rect 554 2623 557 2706
rect 538 2613 557 2616
rect 530 2593 541 2596
rect 578 2593 581 2626
rect 522 2503 525 2526
rect 538 2496 541 2593
rect 530 2493 541 2496
rect 394 2413 421 2416
rect 386 2333 389 2396
rect 386 2303 389 2326
rect 394 2313 397 2413
rect 402 2333 405 2406
rect 410 2393 413 2406
rect 426 2336 429 2406
rect 442 2383 445 2436
rect 450 2423 453 2436
rect 450 2403 453 2416
rect 482 2406 485 2426
rect 478 2403 485 2406
rect 426 2333 445 2336
rect 402 2313 405 2326
rect 378 2213 381 2236
rect 386 2213 389 2226
rect 402 2213 405 2296
rect 290 2193 293 2206
rect 322 2193 325 2206
rect 354 2203 365 2206
rect 362 2193 365 2203
rect 66 2013 69 2026
rect 82 2016 85 2136
rect 74 2013 85 2016
rect 90 2023 117 2026
rect 90 2013 93 2023
rect 122 2016 125 2126
rect 74 1996 77 2013
rect 70 1993 77 1996
rect 70 1896 73 1993
rect 82 1933 85 2006
rect 98 1983 101 2006
rect 106 1943 109 2016
rect 114 2013 125 2016
rect 114 2003 117 2013
rect 82 1903 85 1926
rect 70 1893 77 1896
rect 74 1753 77 1893
rect 90 1813 93 1826
rect 106 1823 109 1926
rect 114 1916 117 1986
rect 130 1983 133 2016
rect 146 2013 149 2026
rect 154 1993 157 2016
rect 162 2003 165 2126
rect 170 2113 173 2136
rect 186 2123 189 2136
rect 122 1923 125 1936
rect 130 1933 133 1956
rect 170 1933 173 1986
rect 178 1933 181 2066
rect 186 2056 189 2116
rect 194 2063 197 2126
rect 186 2053 197 2056
rect 194 2013 197 2053
rect 202 2046 205 2136
rect 226 2133 237 2136
rect 210 2113 213 2126
rect 202 2043 221 2046
rect 202 2023 205 2043
rect 186 1953 189 2006
rect 210 1986 213 2016
rect 218 1993 221 2043
rect 226 2026 229 2126
rect 234 2036 237 2133
rect 266 2123 269 2136
rect 314 2086 317 2136
rect 338 2133 341 2186
rect 386 2123 389 2146
rect 410 2116 413 2326
rect 442 2323 445 2333
rect 418 2303 421 2316
rect 450 2313 453 2326
rect 458 2293 461 2326
rect 466 2313 469 2386
rect 478 2336 481 2403
rect 478 2333 485 2336
rect 418 2223 421 2246
rect 426 2213 429 2226
rect 434 2216 437 2236
rect 442 2223 445 2236
rect 434 2213 453 2216
rect 418 2123 421 2136
rect 426 2133 429 2146
rect 450 2133 453 2196
rect 466 2163 469 2246
rect 474 2203 477 2316
rect 482 2243 485 2333
rect 490 2313 493 2436
rect 530 2433 533 2493
rect 546 2413 549 2426
rect 570 2403 573 2546
rect 586 2523 589 2616
rect 594 2583 597 2816
rect 618 2813 621 2833
rect 602 2713 605 2796
rect 610 2733 613 2806
rect 618 2793 621 2806
rect 626 2803 629 2936
rect 634 2923 637 2946
rect 642 2923 645 2956
rect 650 2923 653 2936
rect 666 2933 669 2946
rect 690 2933 693 2966
rect 746 2936 749 3040
rect 834 2946 837 3040
rect 818 2943 837 2946
rect 658 2846 661 2926
rect 654 2843 661 2846
rect 634 2813 637 2826
rect 634 2793 637 2806
rect 642 2783 645 2816
rect 654 2746 657 2843
rect 610 2696 613 2726
rect 606 2693 613 2696
rect 606 2626 609 2693
rect 618 2633 621 2736
rect 634 2706 637 2746
rect 626 2703 637 2706
rect 650 2743 657 2746
rect 606 2623 613 2626
rect 610 2603 613 2623
rect 618 2553 621 2616
rect 626 2603 629 2703
rect 634 2613 637 2636
rect 650 2623 653 2743
rect 658 2703 661 2736
rect 666 2733 669 2836
rect 674 2726 677 2816
rect 682 2803 685 2926
rect 698 2913 701 2926
rect 714 2896 717 2936
rect 730 2933 749 2936
rect 730 2896 733 2933
rect 738 2913 741 2926
rect 746 2913 749 2926
rect 706 2893 717 2896
rect 722 2893 733 2896
rect 706 2836 709 2893
rect 706 2833 717 2836
rect 690 2813 693 2826
rect 714 2813 717 2833
rect 722 2743 725 2893
rect 730 2823 733 2886
rect 754 2883 757 2916
rect 762 2903 765 2936
rect 770 2913 773 2926
rect 778 2913 781 2926
rect 786 2913 789 2926
rect 794 2923 805 2926
rect 682 2733 693 2736
rect 666 2723 677 2726
rect 666 2713 669 2723
rect 682 2686 685 2726
rect 706 2723 709 2736
rect 682 2683 693 2686
rect 634 2603 653 2606
rect 610 2533 613 2546
rect 626 2533 629 2596
rect 586 2413 589 2426
rect 602 2413 605 2436
rect 610 2403 613 2526
rect 634 2523 637 2603
rect 666 2593 669 2636
rect 690 2613 693 2683
rect 722 2616 725 2696
rect 714 2613 725 2616
rect 642 2496 645 2586
rect 650 2523 653 2536
rect 658 2533 661 2556
rect 634 2493 645 2496
rect 634 2406 637 2493
rect 658 2456 661 2516
rect 666 2513 669 2536
rect 698 2533 701 2606
rect 706 2523 709 2536
rect 730 2533 733 2806
rect 738 2783 741 2816
rect 738 2693 741 2746
rect 714 2513 717 2526
rect 746 2513 749 2826
rect 762 2803 765 2836
rect 754 2723 757 2746
rect 770 2703 773 2826
rect 778 2806 781 2846
rect 818 2843 821 2943
rect 794 2833 805 2836
rect 786 2813 789 2826
rect 794 2813 797 2826
rect 802 2813 805 2833
rect 818 2823 821 2836
rect 826 2806 829 2836
rect 834 2813 837 2926
rect 858 2826 861 3040
rect 890 2913 893 2926
rect 946 2923 949 2946
rect 970 2866 973 2936
rect 986 2913 989 2936
rect 1010 2933 1013 2946
rect 1010 2886 1013 2916
rect 1042 2906 1045 2936
rect 1042 2903 1053 2906
rect 1010 2883 1021 2886
rect 970 2863 981 2866
rect 842 2813 845 2826
rect 858 2823 869 2826
rect 778 2803 789 2806
rect 810 2803 829 2806
rect 786 2723 789 2803
rect 826 2773 829 2803
rect 810 2733 813 2746
rect 866 2736 869 2823
rect 898 2813 901 2826
rect 954 2793 957 2816
rect 834 2733 845 2736
rect 866 2733 877 2736
rect 882 2733 885 2746
rect 754 2626 757 2646
rect 754 2623 761 2626
rect 758 2506 761 2623
rect 770 2593 773 2616
rect 754 2503 761 2506
rect 658 2453 669 2456
rect 634 2403 645 2406
rect 642 2383 645 2403
rect 666 2376 669 2453
rect 714 2433 725 2436
rect 682 2393 685 2416
rect 706 2403 709 2416
rect 658 2373 669 2376
rect 658 2356 661 2373
rect 654 2353 661 2356
rect 498 2323 501 2346
rect 546 2333 557 2336
rect 562 2333 573 2336
rect 514 2223 517 2316
rect 538 2293 541 2316
rect 562 2296 565 2333
rect 570 2313 573 2326
rect 562 2293 573 2296
rect 530 2206 533 2216
rect 482 2193 485 2206
rect 506 2173 509 2206
rect 522 2203 533 2206
rect 562 2193 565 2216
rect 570 2173 573 2293
rect 586 2246 589 2336
rect 610 2323 613 2336
rect 654 2296 657 2353
rect 666 2303 669 2326
rect 674 2313 677 2326
rect 654 2293 661 2296
rect 582 2243 589 2246
rect 582 2196 585 2243
rect 626 2213 629 2226
rect 582 2193 589 2196
rect 458 2133 469 2136
rect 482 2123 501 2126
rect 410 2113 429 2116
rect 314 2083 325 2086
rect 234 2033 253 2036
rect 226 2023 245 2026
rect 210 1983 229 1986
rect 114 1913 125 1916
rect 130 1913 133 1926
rect 98 1813 109 1816
rect 122 1813 125 1913
rect 162 1876 165 1926
rect 162 1873 173 1876
rect 170 1823 173 1873
rect 98 1806 101 1813
rect 82 1803 101 1806
rect 66 1496 69 1716
rect 82 1593 85 1766
rect 106 1723 109 1806
rect 138 1793 141 1806
rect 146 1783 149 1806
rect 114 1706 117 1746
rect 110 1703 117 1706
rect 110 1616 113 1703
rect 110 1613 117 1616
rect 82 1533 85 1586
rect 66 1493 77 1496
rect 74 1346 77 1493
rect 106 1436 109 1596
rect 114 1566 117 1613
rect 122 1583 125 1756
rect 162 1723 165 1796
rect 170 1733 173 1806
rect 178 1793 181 1806
rect 186 1786 189 1926
rect 194 1923 197 1936
rect 202 1926 205 1946
rect 218 1933 221 1946
rect 226 1933 229 1983
rect 234 1943 237 1976
rect 242 1933 245 2023
rect 250 1933 253 2033
rect 258 2003 261 2016
rect 202 1923 213 1926
rect 202 1813 205 1916
rect 210 1803 213 1923
rect 218 1893 221 1926
rect 258 1916 261 1996
rect 266 1983 269 2016
rect 274 1963 277 2006
rect 290 2003 293 2016
rect 314 1996 317 2016
rect 322 2013 325 2083
rect 306 1993 317 1996
rect 290 1976 293 1986
rect 290 1973 301 1976
rect 274 1916 277 1936
rect 250 1913 261 1916
rect 270 1913 277 1916
rect 250 1836 253 1913
rect 250 1833 257 1836
rect 178 1783 189 1786
rect 218 1783 221 1796
rect 178 1733 181 1783
rect 130 1593 133 1616
rect 114 1563 121 1566
rect 118 1506 121 1563
rect 130 1523 133 1546
rect 118 1503 125 1506
rect 102 1433 109 1436
rect 66 1343 77 1346
rect 66 1003 69 1343
rect 82 1203 85 1326
rect 90 1323 93 1406
rect 102 1336 105 1433
rect 122 1426 125 1503
rect 146 1476 149 1616
rect 162 1603 165 1616
rect 178 1613 181 1626
rect 194 1616 197 1766
rect 226 1763 229 1816
rect 242 1783 245 1816
rect 218 1733 221 1756
rect 254 1746 257 1833
rect 270 1826 273 1913
rect 282 1906 285 1926
rect 290 1923 293 1936
rect 298 1923 301 1973
rect 306 1933 309 1993
rect 314 1913 317 1966
rect 282 1903 301 1906
rect 270 1823 277 1826
rect 254 1743 261 1746
rect 202 1713 205 1726
rect 186 1613 197 1616
rect 202 1606 205 1626
rect 170 1536 173 1606
rect 114 1423 125 1426
rect 138 1473 149 1476
rect 154 1533 173 1536
rect 178 1536 181 1606
rect 186 1593 189 1606
rect 194 1603 205 1606
rect 178 1533 189 1536
rect 114 1346 117 1423
rect 138 1406 141 1473
rect 130 1403 141 1406
rect 114 1343 121 1346
rect 98 1333 105 1336
rect 98 1256 101 1333
rect 90 1253 101 1256
rect 90 1196 93 1253
rect 98 1223 101 1246
rect 106 1233 109 1326
rect 118 1256 121 1343
rect 130 1316 133 1403
rect 154 1396 157 1533
rect 162 1413 165 1526
rect 170 1523 173 1533
rect 178 1516 181 1526
rect 170 1513 181 1516
rect 138 1393 157 1396
rect 138 1333 141 1366
rect 146 1343 149 1393
rect 154 1333 157 1346
rect 162 1326 165 1356
rect 170 1346 173 1513
rect 186 1446 189 1533
rect 194 1523 197 1603
rect 202 1533 205 1546
rect 210 1536 213 1606
rect 218 1603 221 1726
rect 242 1723 245 1736
rect 258 1723 261 1743
rect 266 1733 269 1806
rect 274 1803 277 1823
rect 282 1766 285 1896
rect 290 1823 293 1886
rect 298 1793 301 1903
rect 322 1886 325 1946
rect 330 1943 333 1956
rect 338 1933 349 1936
rect 354 1933 357 1946
rect 370 1936 373 2016
rect 386 2003 389 2016
rect 370 1933 381 1936
rect 330 1913 333 1926
rect 314 1883 325 1886
rect 338 1883 341 1933
rect 346 1923 357 1926
rect 282 1763 289 1766
rect 286 1686 289 1763
rect 298 1723 301 1736
rect 306 1723 309 1836
rect 314 1823 317 1883
rect 322 1823 325 1856
rect 322 1813 341 1816
rect 314 1743 317 1806
rect 282 1683 289 1686
rect 226 1603 229 1616
rect 234 1603 237 1626
rect 242 1543 245 1646
rect 282 1643 285 1683
rect 250 1593 253 1606
rect 210 1533 221 1536
rect 226 1533 245 1536
rect 210 1523 221 1526
rect 178 1443 189 1446
rect 178 1353 181 1443
rect 194 1413 197 1426
rect 170 1343 189 1346
rect 170 1333 173 1343
rect 162 1323 173 1326
rect 130 1313 141 1316
rect 114 1253 121 1256
rect 82 1193 93 1196
rect 82 1076 85 1193
rect 114 1176 117 1253
rect 122 1223 125 1236
rect 130 1213 133 1226
rect 110 1173 117 1176
rect 110 1086 113 1173
rect 138 1166 141 1313
rect 146 1206 149 1226
rect 162 1213 165 1266
rect 170 1236 173 1256
rect 178 1243 181 1336
rect 170 1233 181 1236
rect 146 1203 157 1206
rect 106 1083 113 1086
rect 122 1163 141 1166
rect 82 1073 93 1076
rect 90 976 93 1073
rect 82 973 93 976
rect 82 956 85 973
rect 66 953 85 956
rect 106 956 109 1083
rect 106 953 117 956
rect 66 856 69 953
rect 82 933 85 953
rect 82 876 85 926
rect 114 886 117 953
rect 106 883 117 886
rect 82 873 93 876
rect 66 853 77 856
rect 74 796 77 853
rect 66 793 77 796
rect 66 556 69 793
rect 90 776 93 873
rect 82 773 93 776
rect 82 686 85 773
rect 106 756 109 883
rect 106 753 113 756
rect 110 706 113 753
rect 122 716 125 1163
rect 130 1076 133 1126
rect 130 1073 149 1076
rect 138 1013 141 1026
rect 130 983 133 1006
rect 146 1003 149 1073
rect 162 1033 165 1156
rect 170 1113 173 1226
rect 178 1153 181 1233
rect 186 1223 189 1326
rect 194 1313 197 1326
rect 178 1123 181 1146
rect 186 1116 189 1216
rect 194 1213 197 1236
rect 194 1123 197 1166
rect 178 1113 189 1116
rect 154 1013 165 1016
rect 170 1006 173 1016
rect 130 923 133 946
rect 138 813 141 826
rect 130 783 133 806
rect 146 766 149 806
rect 130 763 149 766
rect 130 723 133 763
rect 154 746 157 1006
rect 162 1003 173 1006
rect 162 923 165 996
rect 170 906 173 1003
rect 178 986 181 1113
rect 202 1103 205 1416
rect 210 1346 213 1523
rect 234 1516 237 1533
rect 230 1513 237 1516
rect 230 1436 233 1513
rect 230 1433 237 1436
rect 218 1376 221 1426
rect 226 1403 229 1416
rect 218 1373 229 1376
rect 210 1343 221 1346
rect 210 1223 213 1336
rect 218 1253 221 1343
rect 226 1333 229 1373
rect 234 1313 237 1433
rect 242 1413 245 1516
rect 250 1333 253 1406
rect 258 1333 261 1636
rect 266 1603 269 1616
rect 282 1613 285 1626
rect 306 1613 309 1716
rect 314 1706 317 1736
rect 322 1713 325 1726
rect 338 1723 341 1813
rect 346 1733 349 1846
rect 354 1813 357 1923
rect 378 1913 381 1933
rect 378 1883 381 1906
rect 386 1856 389 1926
rect 386 1853 397 1856
rect 354 1793 357 1806
rect 378 1803 381 1826
rect 394 1823 397 1853
rect 386 1796 389 1816
rect 402 1803 405 1946
rect 410 1933 413 2016
rect 426 1876 429 2026
rect 466 2006 469 2016
rect 474 2013 477 2026
rect 466 2003 485 2006
rect 434 1913 437 1946
rect 442 1903 445 1946
rect 482 1936 485 2003
rect 490 1943 493 2006
rect 450 1923 453 1936
rect 474 1926 477 1936
rect 482 1933 493 1936
rect 498 1933 501 2123
rect 418 1873 429 1876
rect 410 1813 413 1826
rect 418 1823 421 1873
rect 426 1813 429 1826
rect 378 1793 389 1796
rect 314 1703 325 1706
rect 354 1703 357 1726
rect 322 1613 325 1703
rect 274 1553 277 1606
rect 290 1546 293 1606
rect 298 1593 301 1606
rect 314 1593 317 1606
rect 274 1543 293 1546
rect 266 1506 269 1526
rect 298 1523 301 1536
rect 266 1503 277 1506
rect 274 1446 277 1503
rect 266 1443 277 1446
rect 306 1446 309 1536
rect 314 1533 317 1546
rect 306 1443 317 1446
rect 218 1223 221 1246
rect 226 1216 229 1236
rect 210 1213 229 1216
rect 234 1206 237 1276
rect 242 1213 245 1326
rect 250 1313 253 1326
rect 250 1223 253 1306
rect 226 1203 237 1206
rect 218 1133 221 1146
rect 210 1113 213 1126
rect 226 1116 229 1203
rect 222 1113 229 1116
rect 186 993 189 1006
rect 178 983 197 986
rect 178 926 181 976
rect 186 933 189 946
rect 178 923 189 926
rect 166 903 173 906
rect 166 826 169 903
rect 166 823 173 826
rect 170 803 173 823
rect 178 796 181 916
rect 186 813 189 923
rect 194 906 197 983
rect 202 973 205 1036
rect 210 933 213 1026
rect 222 976 225 1113
rect 234 983 237 1126
rect 222 973 229 976
rect 194 903 205 906
rect 202 856 205 903
rect 194 853 205 856
rect 194 813 197 853
rect 218 836 221 946
rect 226 913 229 973
rect 242 923 245 1206
rect 258 1163 261 1326
rect 266 1303 269 1443
rect 274 1283 277 1416
rect 290 1413 293 1426
rect 266 1216 269 1236
rect 274 1223 277 1236
rect 282 1223 285 1376
rect 290 1313 293 1406
rect 290 1246 293 1286
rect 298 1253 301 1316
rect 306 1273 309 1406
rect 314 1373 317 1443
rect 322 1403 325 1606
rect 330 1543 333 1606
rect 346 1556 349 1606
rect 362 1563 365 1736
rect 378 1723 381 1793
rect 386 1733 397 1736
rect 418 1733 421 1806
rect 386 1633 389 1733
rect 394 1723 413 1726
rect 434 1723 437 1816
rect 442 1813 445 1826
rect 466 1823 469 1926
rect 474 1923 485 1926
rect 474 1903 477 1916
rect 474 1823 477 1856
rect 482 1843 485 1923
rect 450 1813 477 1816
rect 442 1793 445 1806
rect 450 1733 453 1813
rect 474 1776 477 1806
rect 482 1783 485 1806
rect 490 1793 493 1933
rect 506 1906 509 2026
rect 522 2003 525 2126
rect 538 2013 541 2026
rect 562 2023 565 2136
rect 586 2133 589 2193
rect 610 2143 613 2206
rect 626 2123 629 2206
rect 650 2173 653 2206
rect 658 2123 661 2293
rect 682 2273 685 2326
rect 690 2313 693 2336
rect 698 2333 701 2346
rect 682 2213 685 2226
rect 698 2223 701 2266
rect 706 2243 709 2386
rect 722 2343 725 2426
rect 730 2423 733 2436
rect 738 2413 741 2426
rect 754 2386 757 2503
rect 762 2393 765 2406
rect 770 2403 773 2526
rect 754 2383 765 2386
rect 722 2266 725 2336
rect 714 2263 725 2266
rect 666 2123 669 2206
rect 674 2133 677 2206
rect 698 2203 701 2216
rect 714 2173 717 2263
rect 738 2176 741 2216
rect 746 2213 749 2326
rect 754 2206 757 2246
rect 722 2173 741 2176
rect 746 2203 757 2206
rect 682 2123 701 2126
rect 706 2113 709 2166
rect 722 2133 725 2173
rect 738 2133 741 2146
rect 746 2133 749 2203
rect 762 2176 765 2383
rect 778 2366 781 2416
rect 786 2403 789 2426
rect 794 2396 797 2726
rect 810 2626 813 2726
rect 834 2636 837 2733
rect 842 2703 845 2726
rect 850 2713 853 2726
rect 858 2663 861 2726
rect 866 2703 869 2726
rect 834 2633 845 2636
rect 810 2623 837 2626
rect 810 2523 813 2623
rect 818 2603 821 2616
rect 834 2593 837 2606
rect 842 2533 845 2633
rect 858 2583 861 2616
rect 874 2613 877 2733
rect 890 2723 893 2776
rect 978 2756 981 2863
rect 1018 2836 1021 2883
rect 994 2803 997 2826
rect 970 2753 981 2756
rect 946 2723 949 2736
rect 970 2676 973 2753
rect 986 2733 989 2776
rect 1002 2723 1005 2816
rect 1010 2813 1013 2836
rect 1018 2833 1037 2836
rect 1018 2823 1021 2833
rect 1026 2813 1029 2826
rect 1010 2723 1013 2746
rect 1018 2733 1021 2806
rect 1034 2766 1037 2833
rect 1050 2816 1053 2903
rect 1058 2823 1061 2836
rect 1042 2783 1045 2816
rect 1050 2813 1061 2816
rect 1050 2786 1053 2813
rect 1058 2793 1061 2806
rect 1066 2803 1069 2946
rect 1082 2803 1085 2816
rect 1050 2783 1057 2786
rect 1026 2763 1037 2766
rect 1026 2716 1029 2763
rect 1002 2713 1029 2716
rect 1054 2716 1057 2783
rect 1066 2723 1069 2746
rect 1054 2713 1061 2716
rect 1026 2686 1029 2713
rect 1026 2683 1045 2686
rect 970 2673 981 2676
rect 970 2623 973 2666
rect 866 2543 869 2606
rect 930 2593 933 2616
rect 954 2573 957 2606
rect 970 2593 973 2606
rect 978 2586 981 2673
rect 1042 2666 1045 2683
rect 1042 2663 1049 2666
rect 962 2583 981 2586
rect 834 2433 837 2526
rect 842 2503 845 2516
rect 850 2503 853 2516
rect 858 2486 861 2526
rect 874 2523 885 2526
rect 858 2483 869 2486
rect 826 2423 837 2426
rect 794 2393 801 2396
rect 778 2363 789 2366
rect 762 2173 773 2176
rect 754 2133 765 2136
rect 730 2123 741 2126
rect 514 1933 517 1956
rect 522 1933 533 1936
rect 538 1933 541 2006
rect 546 1953 549 2006
rect 514 1913 517 1926
rect 498 1903 509 1906
rect 498 1823 501 1903
rect 498 1783 501 1816
rect 506 1793 509 1836
rect 522 1813 525 1926
rect 530 1833 533 1926
rect 546 1893 549 1926
rect 554 1903 557 1966
rect 562 1943 565 2016
rect 586 1963 589 2016
rect 562 1923 565 1936
rect 578 1893 581 1926
rect 474 1773 493 1776
rect 466 1733 477 1736
rect 482 1723 485 1736
rect 490 1723 493 1773
rect 538 1753 541 1806
rect 394 1703 397 1716
rect 474 1703 477 1716
rect 386 1593 389 1616
rect 434 1593 437 1606
rect 458 1566 461 1676
rect 498 1613 501 1736
rect 514 1726 517 1736
rect 522 1733 525 1746
rect 562 1733 565 1756
rect 578 1733 581 1816
rect 586 1813 589 1936
rect 618 1926 621 1956
rect 626 1933 629 1946
rect 634 1933 637 2016
rect 666 2013 669 2026
rect 610 1913 613 1926
rect 618 1923 629 1926
rect 650 1923 653 2006
rect 658 1933 661 1976
rect 674 1973 677 2016
rect 682 1953 685 2006
rect 690 2003 693 2026
rect 698 2003 701 2016
rect 666 1923 669 1936
rect 682 1926 685 1946
rect 674 1923 685 1926
rect 626 1853 629 1923
rect 634 1913 645 1916
rect 634 1826 637 1913
rect 690 1873 693 1936
rect 698 1933 717 1936
rect 698 1913 701 1933
rect 706 1923 733 1926
rect 738 1923 741 2116
rect 762 2113 765 2126
rect 770 2083 773 2173
rect 778 2126 781 2246
rect 786 2183 789 2363
rect 798 2266 801 2393
rect 794 2263 801 2266
rect 794 2243 797 2263
rect 794 2143 797 2216
rect 802 2213 805 2226
rect 810 2213 813 2346
rect 818 2323 821 2406
rect 826 2323 829 2423
rect 834 2413 853 2416
rect 826 2193 829 2226
rect 834 2213 837 2413
rect 802 2143 805 2166
rect 842 2156 845 2236
rect 826 2153 845 2156
rect 778 2123 789 2126
rect 786 2076 789 2123
rect 810 2093 813 2116
rect 818 2103 821 2136
rect 826 2123 829 2153
rect 842 2133 845 2146
rect 834 2086 837 2126
rect 842 2113 845 2126
rect 850 2123 853 2336
rect 858 2323 861 2436
rect 866 2413 869 2483
rect 874 2423 877 2516
rect 898 2423 909 2426
rect 922 2423 925 2436
rect 938 2423 941 2526
rect 962 2463 965 2583
rect 978 2533 981 2546
rect 994 2533 997 2606
rect 1002 2603 1005 2616
rect 1018 2603 1021 2616
rect 1046 2596 1049 2663
rect 1042 2593 1049 2596
rect 1042 2573 1045 2593
rect 1010 2533 1013 2546
rect 866 2403 877 2406
rect 890 2383 893 2416
rect 898 2413 917 2416
rect 898 2403 901 2413
rect 938 2366 941 2406
rect 930 2363 941 2366
rect 866 2333 869 2346
rect 866 2323 885 2326
rect 890 2303 893 2336
rect 906 2323 917 2326
rect 866 2206 869 2236
rect 882 2213 885 2226
rect 898 2213 901 2316
rect 930 2313 933 2363
rect 906 2213 909 2226
rect 922 2223 925 2236
rect 866 2203 885 2206
rect 898 2203 909 2206
rect 922 2203 925 2216
rect 938 2213 941 2346
rect 946 2213 949 2326
rect 954 2316 957 2396
rect 978 2393 981 2406
rect 986 2403 989 2416
rect 994 2413 997 2526
rect 1018 2406 1021 2536
rect 1026 2413 1029 2426
rect 1010 2326 1013 2406
rect 1018 2403 1029 2406
rect 1050 2403 1053 2526
rect 1058 2523 1061 2713
rect 1066 2593 1069 2616
rect 1090 2546 1093 2846
rect 1106 2813 1109 2836
rect 1106 2636 1109 2806
rect 1114 2723 1117 2916
rect 1122 2856 1125 2926
rect 1122 2853 1133 2856
rect 1130 2803 1133 2853
rect 1146 2843 1149 2936
rect 1162 2933 1165 3040
rect 1234 2966 1237 3040
rect 1230 2963 1237 2966
rect 1170 2943 1181 2946
rect 1162 2913 1165 2926
rect 1138 2823 1165 2826
rect 1138 2803 1141 2816
rect 1162 2813 1165 2823
rect 1178 2813 1181 2936
rect 1194 2933 1213 2936
rect 1194 2833 1197 2933
rect 1202 2916 1205 2926
rect 1210 2923 1213 2933
rect 1218 2916 1221 2926
rect 1202 2913 1221 2916
rect 1230 2886 1233 2963
rect 1298 2943 1301 3040
rect 1378 2966 1381 3040
rect 1458 3026 1461 3040
rect 1450 3023 1461 3026
rect 1450 2976 1453 3023
rect 1450 2973 1461 2976
rect 1370 2963 1381 2966
rect 1230 2883 1237 2886
rect 1194 2813 1197 2826
rect 1154 2793 1157 2806
rect 1170 2773 1173 2806
rect 1178 2793 1181 2806
rect 1202 2796 1205 2826
rect 1210 2813 1213 2846
rect 1218 2813 1221 2836
rect 1234 2823 1237 2883
rect 1226 2803 1229 2816
rect 1202 2793 1221 2796
rect 1122 2706 1125 2736
rect 1130 2733 1133 2746
rect 1138 2723 1141 2736
rect 1146 2723 1149 2736
rect 1186 2733 1189 2756
rect 1154 2716 1157 2726
rect 1130 2713 1157 2716
rect 1162 2716 1165 2726
rect 1162 2713 1169 2716
rect 1122 2703 1133 2706
rect 1082 2543 1093 2546
rect 1098 2633 1109 2636
rect 1074 2503 1077 2526
rect 1082 2436 1085 2543
rect 1090 2523 1093 2536
rect 1098 2523 1101 2633
rect 1106 2623 1125 2626
rect 1106 2613 1109 2623
rect 1114 2603 1117 2616
rect 1122 2613 1125 2623
rect 1130 2596 1133 2703
rect 1166 2636 1169 2713
rect 1138 2603 1141 2616
rect 1146 2606 1149 2626
rect 1154 2616 1157 2636
rect 1166 2633 1173 2636
rect 1154 2613 1165 2616
rect 1146 2603 1157 2606
rect 1130 2593 1141 2596
rect 1162 2546 1165 2613
rect 1170 2603 1173 2633
rect 1178 2613 1181 2726
rect 1194 2696 1197 2736
rect 1186 2693 1197 2696
rect 1186 2613 1189 2693
rect 1202 2623 1205 2726
rect 1218 2723 1221 2793
rect 1234 2763 1237 2816
rect 1242 2813 1253 2816
rect 1258 2786 1261 2826
rect 1266 2803 1269 2926
rect 1298 2923 1301 2936
rect 1274 2826 1277 2846
rect 1274 2823 1281 2826
rect 1242 2783 1261 2786
rect 1234 2733 1237 2746
rect 1242 2723 1245 2783
rect 1250 2733 1253 2766
rect 1258 2723 1261 2776
rect 1266 2643 1269 2756
rect 1278 2746 1281 2823
rect 1290 2813 1293 2846
rect 1290 2793 1293 2806
rect 1298 2803 1309 2806
rect 1298 2783 1301 2803
rect 1274 2743 1281 2746
rect 1274 2653 1277 2743
rect 1290 2733 1301 2736
rect 1282 2663 1285 2726
rect 1314 2723 1317 2946
rect 1330 2923 1333 2936
rect 1322 2793 1325 2806
rect 1330 2783 1333 2826
rect 1338 2793 1341 2846
rect 1346 2786 1349 2806
rect 1338 2783 1349 2786
rect 1338 2743 1341 2783
rect 1194 2613 1205 2616
rect 1218 2613 1221 2636
rect 1266 2623 1269 2636
rect 1194 2606 1197 2613
rect 1178 2603 1197 2606
rect 1202 2593 1205 2606
rect 1226 2593 1229 2606
rect 1234 2583 1237 2606
rect 1242 2603 1245 2616
rect 1258 2593 1261 2606
rect 1266 2583 1269 2616
rect 1290 2606 1293 2616
rect 1274 2603 1293 2606
rect 1298 2603 1301 2646
rect 1306 2613 1309 2636
rect 1154 2533 1157 2546
rect 1162 2543 1173 2546
rect 1130 2513 1133 2526
rect 1162 2503 1165 2536
rect 1082 2433 1101 2436
rect 1026 2393 1029 2403
rect 1034 2356 1037 2396
rect 1026 2353 1037 2356
rect 1018 2333 1021 2346
rect 1026 2333 1029 2353
rect 962 2323 981 2326
rect 954 2313 973 2316
rect 978 2303 981 2323
rect 986 2233 989 2326
rect 994 2313 997 2326
rect 1010 2323 1021 2326
rect 1026 2323 1045 2326
rect 1058 2323 1061 2336
rect 1002 2303 1005 2316
rect 1018 2313 1021 2323
rect 1066 2286 1069 2346
rect 1074 2323 1077 2416
rect 1082 2336 1085 2356
rect 1098 2353 1101 2433
rect 1146 2393 1149 2416
rect 1170 2366 1173 2543
rect 1178 2496 1181 2526
rect 1194 2523 1197 2576
rect 1202 2506 1205 2546
rect 1218 2533 1229 2536
rect 1198 2503 1205 2506
rect 1178 2493 1189 2496
rect 1186 2396 1189 2493
rect 1198 2406 1201 2503
rect 1210 2423 1213 2526
rect 1226 2523 1245 2526
rect 1266 2523 1269 2536
rect 1274 2523 1277 2603
rect 1306 2593 1309 2606
rect 1314 2583 1317 2606
rect 1322 2556 1325 2736
rect 1354 2733 1357 2926
rect 1370 2886 1373 2963
rect 1370 2883 1381 2886
rect 1362 2813 1365 2836
rect 1370 2796 1373 2816
rect 1378 2806 1381 2883
rect 1410 2833 1413 2926
rect 1426 2876 1429 2936
rect 1418 2873 1429 2876
rect 1378 2803 1389 2806
rect 1370 2793 1381 2796
rect 1338 2623 1341 2666
rect 1370 2646 1373 2786
rect 1378 2733 1381 2793
rect 1386 2693 1389 2803
rect 1418 2766 1421 2873
rect 1458 2863 1461 2973
rect 1474 2966 1477 3040
rect 1474 2963 1493 2966
rect 1474 2923 1477 2946
rect 1490 2886 1493 2963
rect 1498 2926 1501 3040
rect 1498 2923 1509 2926
rect 1486 2883 1493 2886
rect 1486 2826 1489 2883
rect 1482 2823 1489 2826
rect 1466 2803 1469 2816
rect 1402 2763 1421 2766
rect 1370 2643 1381 2646
rect 1338 2556 1341 2606
rect 1346 2603 1349 2626
rect 1354 2613 1357 2636
rect 1378 2613 1381 2643
rect 1314 2553 1325 2556
rect 1330 2553 1341 2556
rect 1226 2416 1229 2516
rect 1210 2413 1229 2416
rect 1198 2403 1205 2406
rect 1178 2393 1189 2396
rect 1178 2373 1181 2393
rect 1202 2386 1205 2403
rect 1210 2393 1213 2406
rect 1202 2383 1221 2386
rect 1162 2363 1173 2366
rect 1082 2333 1093 2336
rect 1074 2293 1077 2316
rect 1066 2283 1077 2286
rect 1002 2233 1021 2236
rect 978 2223 989 2226
rect 986 2216 989 2223
rect 1002 2216 1005 2233
rect 858 2133 861 2156
rect 866 2123 869 2186
rect 906 2163 909 2203
rect 946 2193 949 2206
rect 970 2203 973 2216
rect 978 2203 981 2216
rect 986 2213 1005 2216
rect 1010 2213 1013 2226
rect 1018 2213 1021 2233
rect 834 2083 845 2086
rect 778 2073 789 2076
rect 778 2033 781 2073
rect 746 1996 749 2016
rect 754 2003 757 2016
rect 746 1993 773 1996
rect 770 1983 773 1993
rect 610 1823 637 1826
rect 506 1693 509 1726
rect 514 1723 525 1726
rect 338 1553 349 1556
rect 338 1523 341 1553
rect 330 1413 333 1436
rect 346 1426 349 1536
rect 354 1513 357 1526
rect 362 1523 365 1546
rect 370 1513 373 1536
rect 346 1423 373 1426
rect 314 1266 317 1326
rect 322 1313 325 1386
rect 306 1263 317 1266
rect 290 1243 301 1246
rect 266 1213 285 1216
rect 298 1213 301 1243
rect 306 1203 309 1263
rect 314 1203 317 1226
rect 250 1126 253 1146
rect 282 1143 293 1146
rect 250 1123 261 1126
rect 290 1123 293 1143
rect 258 1046 261 1123
rect 298 1103 301 1136
rect 306 1113 309 1136
rect 322 1133 325 1246
rect 330 1223 333 1406
rect 346 1393 349 1423
rect 354 1413 373 1416
rect 354 1383 357 1406
rect 354 1336 357 1346
rect 338 1313 341 1336
rect 354 1333 365 1336
rect 370 1333 373 1413
rect 338 1216 341 1226
rect 346 1223 349 1246
rect 354 1223 357 1326
rect 362 1323 365 1333
rect 370 1313 373 1326
rect 378 1323 381 1536
rect 386 1523 389 1536
rect 394 1436 397 1566
rect 442 1563 461 1566
rect 418 1513 421 1546
rect 442 1486 445 1563
rect 466 1523 469 1556
rect 514 1523 517 1536
rect 538 1533 541 1626
rect 546 1603 549 1726
rect 554 1603 557 1666
rect 570 1643 573 1726
rect 586 1616 589 1806
rect 610 1636 613 1823
rect 618 1733 621 1816
rect 626 1753 629 1806
rect 634 1763 637 1816
rect 642 1793 645 1806
rect 650 1803 653 1816
rect 658 1743 661 1806
rect 674 1783 677 1806
rect 698 1793 701 1816
rect 698 1746 701 1786
rect 682 1743 701 1746
rect 610 1633 617 1636
rect 570 1613 589 1616
rect 602 1613 605 1626
rect 562 1543 565 1606
rect 578 1593 581 1606
rect 554 1533 573 1536
rect 562 1513 565 1526
rect 442 1483 453 1486
rect 386 1433 397 1436
rect 410 1433 421 1436
rect 386 1356 389 1433
rect 410 1426 413 1433
rect 394 1423 413 1426
rect 426 1423 429 1436
rect 394 1413 397 1423
rect 386 1353 397 1356
rect 386 1333 389 1346
rect 394 1236 397 1353
rect 402 1343 405 1416
rect 410 1403 413 1423
rect 426 1413 437 1416
rect 402 1306 405 1326
rect 410 1313 413 1326
rect 402 1303 413 1306
rect 418 1293 421 1326
rect 426 1306 429 1396
rect 434 1333 445 1336
rect 434 1313 437 1333
rect 426 1303 437 1306
rect 362 1216 365 1226
rect 330 1213 341 1216
rect 346 1213 357 1216
rect 362 1213 373 1216
rect 378 1206 381 1236
rect 370 1203 381 1206
rect 386 1233 397 1236
rect 410 1233 413 1256
rect 418 1233 421 1246
rect 386 1196 389 1233
rect 394 1213 397 1226
rect 378 1193 389 1196
rect 394 1193 397 1206
rect 250 1043 261 1046
rect 250 1013 253 1043
rect 250 983 253 996
rect 258 973 261 1006
rect 266 983 269 1006
rect 274 933 277 1006
rect 282 993 285 1016
rect 290 996 293 1046
rect 314 1016 317 1126
rect 338 1123 341 1136
rect 370 1123 373 1136
rect 306 1013 317 1016
rect 338 1013 341 1026
rect 346 1006 349 1106
rect 378 1043 381 1193
rect 402 1186 405 1226
rect 418 1223 429 1226
rect 386 1183 405 1186
rect 386 1123 389 1183
rect 394 1133 397 1146
rect 410 1133 413 1216
rect 434 1213 437 1303
rect 442 1253 445 1326
rect 450 1246 453 1483
rect 458 1286 461 1336
rect 466 1293 469 1326
rect 458 1283 469 1286
rect 442 1243 453 1246
rect 442 1203 445 1243
rect 450 1223 453 1236
rect 370 1013 373 1036
rect 386 1026 389 1116
rect 410 1113 413 1126
rect 418 1083 421 1126
rect 450 1123 453 1146
rect 466 1133 469 1283
rect 474 1233 477 1436
rect 506 1416 509 1426
rect 506 1413 525 1416
rect 498 1336 501 1406
rect 522 1403 525 1413
rect 490 1333 501 1336
rect 482 1303 485 1316
rect 490 1263 493 1333
rect 498 1313 501 1326
rect 506 1313 509 1326
rect 522 1296 525 1336
rect 530 1323 533 1426
rect 538 1413 557 1416
rect 554 1326 557 1336
rect 562 1333 565 1406
rect 570 1403 573 1416
rect 586 1413 589 1606
rect 614 1586 617 1633
rect 626 1593 629 1606
rect 634 1593 637 1606
rect 650 1596 653 1726
rect 682 1713 685 1726
rect 698 1716 701 1736
rect 706 1723 709 1746
rect 694 1713 701 1716
rect 642 1593 653 1596
rect 614 1583 633 1586
rect 610 1533 613 1556
rect 602 1456 605 1526
rect 598 1453 605 1456
rect 578 1393 581 1406
rect 598 1366 601 1453
rect 618 1413 621 1546
rect 630 1506 633 1583
rect 642 1513 645 1593
rect 630 1503 637 1506
rect 598 1363 605 1366
rect 586 1333 589 1356
rect 602 1333 605 1363
rect 538 1313 541 1326
rect 546 1323 557 1326
rect 546 1306 549 1323
rect 562 1316 565 1326
rect 562 1313 573 1316
rect 546 1303 565 1306
rect 522 1293 533 1296
rect 482 1203 485 1256
rect 490 1213 493 1226
rect 498 1223 509 1226
rect 498 1103 501 1136
rect 514 1133 517 1216
rect 522 1123 525 1206
rect 530 1203 533 1293
rect 554 1213 557 1296
rect 450 1043 469 1046
rect 378 1023 389 1026
rect 402 1023 413 1026
rect 418 1023 421 1036
rect 426 1023 429 1036
rect 450 1023 453 1043
rect 290 993 301 996
rect 314 993 317 1006
rect 282 933 285 976
rect 298 926 301 993
rect 322 983 325 1006
rect 330 1003 349 1006
rect 202 833 221 836
rect 150 743 157 746
rect 162 793 181 796
rect 186 793 189 806
rect 122 713 133 716
rect 110 703 117 706
rect 82 683 93 686
rect 90 573 93 683
rect 114 646 117 703
rect 114 643 121 646
rect 118 596 121 643
rect 114 593 121 596
rect 66 553 85 556
rect 82 176 85 553
rect 114 513 117 593
rect 122 496 125 536
rect 114 493 125 496
rect 114 436 117 493
rect 114 433 125 436
rect 122 403 125 433
rect 130 373 133 713
rect 150 666 153 743
rect 162 676 165 793
rect 170 713 173 726
rect 178 723 181 786
rect 194 736 197 806
rect 202 783 205 833
rect 218 763 221 806
rect 242 793 245 816
rect 250 773 253 926
rect 290 923 301 926
rect 290 826 293 923
rect 314 913 317 926
rect 322 893 325 926
rect 330 903 333 1003
rect 338 923 341 996
rect 362 993 365 1006
rect 346 846 349 936
rect 338 843 349 846
rect 286 823 293 826
rect 194 733 201 736
rect 266 733 269 766
rect 162 673 169 676
rect 150 663 157 666
rect 138 576 141 616
rect 138 573 149 576
rect 138 476 141 536
rect 146 533 149 573
rect 154 533 157 663
rect 166 606 169 673
rect 186 626 189 726
rect 198 636 201 733
rect 286 726 289 823
rect 298 813 325 816
rect 298 733 301 813
rect 330 803 333 826
rect 306 773 309 796
rect 242 636 245 726
rect 286 723 293 726
rect 314 723 317 786
rect 330 743 333 756
rect 338 733 341 843
rect 354 836 357 986
rect 362 923 365 936
rect 346 833 357 836
rect 346 803 349 833
rect 354 783 357 816
rect 362 803 365 916
rect 362 733 365 776
rect 370 733 373 976
rect 378 966 381 1023
rect 386 1003 389 1016
rect 394 993 397 1006
rect 402 983 405 1023
rect 410 1013 421 1016
rect 426 1006 429 1016
rect 458 1013 461 1036
rect 426 1003 453 1006
rect 378 963 389 966
rect 378 913 381 926
rect 386 923 389 963
rect 410 923 413 936
rect 378 793 381 816
rect 386 803 389 916
rect 394 896 397 916
rect 394 893 405 896
rect 394 813 397 826
rect 402 823 405 893
rect 410 823 413 836
rect 386 736 389 746
rect 386 733 397 736
rect 338 723 357 726
rect 290 703 293 723
rect 338 713 341 723
rect 386 713 389 726
rect 394 723 397 733
rect 402 706 405 786
rect 198 633 205 636
rect 242 633 253 636
rect 178 613 181 626
rect 186 623 197 626
rect 162 603 169 606
rect 162 583 165 603
rect 162 533 165 546
rect 186 543 189 616
rect 194 593 197 623
rect 138 473 149 476
rect 138 366 141 406
rect 130 363 141 366
rect 130 323 133 363
rect 146 323 149 473
rect 154 413 157 526
rect 154 393 157 406
rect 162 403 165 526
rect 170 513 173 536
rect 170 366 173 476
rect 202 473 205 633
rect 226 603 229 616
rect 234 613 237 626
rect 250 616 253 633
rect 250 613 257 616
rect 234 596 237 606
rect 218 593 237 596
rect 186 413 189 426
rect 154 363 173 366
rect 154 306 157 363
rect 178 343 181 406
rect 194 393 197 416
rect 210 393 213 406
rect 162 323 165 336
rect 178 313 181 336
rect 202 323 205 346
rect 210 326 213 376
rect 218 333 221 406
rect 234 393 237 416
rect 242 373 245 586
rect 254 556 257 613
rect 250 553 257 556
rect 250 533 253 553
rect 266 533 269 616
rect 258 513 261 526
rect 274 523 277 626
rect 298 616 301 626
rect 282 593 285 616
rect 290 613 301 616
rect 298 593 301 606
rect 314 603 317 616
rect 338 606 341 706
rect 402 703 413 706
rect 418 693 421 926
rect 426 923 429 1003
rect 434 846 437 986
rect 466 936 469 1043
rect 474 1033 485 1036
rect 474 1013 477 1033
rect 482 1013 485 1026
rect 466 933 473 936
rect 458 913 461 926
rect 442 893 445 906
rect 470 886 473 933
rect 482 893 485 916
rect 490 913 493 1016
rect 506 936 509 1026
rect 514 1003 517 1086
rect 522 1003 525 1116
rect 530 1033 533 1136
rect 538 1123 541 1136
rect 546 1133 549 1156
rect 562 1126 565 1303
rect 570 1223 573 1313
rect 578 1273 581 1326
rect 594 1213 597 1286
rect 578 1153 581 1206
rect 546 1113 549 1126
rect 554 1123 565 1126
rect 554 1113 557 1123
rect 538 993 541 1106
rect 562 1013 565 1036
rect 578 1026 581 1146
rect 602 1123 605 1326
rect 626 1323 629 1336
rect 634 1323 637 1503
rect 666 1453 669 1616
rect 674 1573 677 1606
rect 682 1533 685 1636
rect 694 1626 697 1713
rect 694 1623 701 1626
rect 698 1583 701 1623
rect 706 1533 709 1706
rect 714 1653 717 1923
rect 722 1713 725 1746
rect 714 1603 717 1616
rect 722 1596 725 1606
rect 730 1603 733 1736
rect 738 1703 741 1826
rect 762 1723 765 1816
rect 770 1783 773 1816
rect 786 1803 789 1966
rect 794 1923 797 1946
rect 818 1933 821 2036
rect 842 2013 845 2083
rect 834 1956 837 2006
rect 850 1993 853 2006
rect 834 1953 845 1956
rect 834 1933 837 1946
rect 842 1933 845 1953
rect 850 1933 853 1956
rect 858 1913 861 1926
rect 866 1853 869 2096
rect 874 2073 877 2136
rect 874 1913 877 2006
rect 882 2003 885 2136
rect 898 2116 901 2136
rect 954 2133 957 2156
rect 978 2133 981 2166
rect 890 2113 901 2116
rect 906 2113 909 2126
rect 898 2013 901 2106
rect 922 2056 925 2126
rect 962 2096 965 2116
rect 954 2093 965 2096
rect 922 2053 933 2056
rect 882 1923 885 1986
rect 890 1953 893 2006
rect 770 1703 773 1736
rect 778 1723 781 1746
rect 794 1733 797 1776
rect 818 1773 821 1836
rect 866 1823 877 1826
rect 882 1816 885 1916
rect 898 1913 901 2006
rect 922 1993 925 2006
rect 930 1993 933 2053
rect 954 2046 957 2093
rect 954 2043 965 2046
rect 954 2013 957 2026
rect 930 1933 933 1956
rect 938 1923 941 1936
rect 946 1933 949 1946
rect 954 1883 957 2006
rect 962 1986 965 2043
rect 970 2013 973 2116
rect 978 2093 981 2126
rect 986 2113 989 2126
rect 994 2103 997 2126
rect 1002 2113 1005 2213
rect 1026 2206 1029 2236
rect 1050 2213 1053 2226
rect 1058 2223 1061 2236
rect 1066 2206 1069 2236
rect 1074 2213 1077 2283
rect 1090 2256 1093 2333
rect 1106 2283 1109 2326
rect 1114 2313 1117 2336
rect 1122 2303 1125 2326
rect 1162 2276 1165 2363
rect 1202 2333 1205 2356
rect 1162 2273 1173 2276
rect 1082 2253 1093 2256
rect 1010 2203 1029 2206
rect 1050 2203 1069 2206
rect 1026 2193 1029 2203
rect 1018 2066 1021 2156
rect 1082 2153 1085 2253
rect 1090 2233 1101 2236
rect 1098 2226 1101 2233
rect 1090 2213 1093 2226
rect 1098 2223 1109 2226
rect 1106 2163 1109 2223
rect 1114 2183 1117 2216
rect 1122 2213 1125 2226
rect 1162 2213 1165 2256
rect 1138 2193 1141 2206
rect 1042 2123 1045 2146
rect 1002 2063 1021 2066
rect 978 1993 981 2006
rect 986 1993 989 2006
rect 1002 2003 1005 2063
rect 1098 2036 1101 2126
rect 1106 2103 1109 2116
rect 1114 2093 1117 2126
rect 1122 2103 1125 2126
rect 1138 2123 1141 2166
rect 1146 2116 1149 2136
rect 1130 2113 1149 2116
rect 1154 2103 1157 2136
rect 1170 2043 1173 2273
rect 1178 2213 1181 2326
rect 1218 2313 1221 2383
rect 1226 2323 1229 2336
rect 1234 2323 1237 2406
rect 1242 2393 1245 2523
rect 1314 2513 1317 2553
rect 1322 2496 1325 2546
rect 1330 2523 1333 2553
rect 1318 2493 1325 2496
rect 1266 2406 1269 2436
rect 1274 2413 1301 2416
rect 1266 2403 1285 2406
rect 1242 2336 1245 2376
rect 1242 2333 1253 2336
rect 1218 2223 1229 2226
rect 1194 2193 1197 2206
rect 1202 2193 1205 2216
rect 1218 2206 1221 2223
rect 1210 2203 1221 2206
rect 1226 2193 1229 2216
rect 1242 2203 1245 2326
rect 1250 2293 1253 2333
rect 1258 2323 1261 2386
rect 1298 2383 1301 2413
rect 1306 2373 1309 2446
rect 1318 2426 1321 2493
rect 1318 2423 1325 2426
rect 1322 2403 1325 2423
rect 1330 2413 1333 2516
rect 1354 2453 1357 2556
rect 1378 2543 1381 2606
rect 1378 2516 1381 2536
rect 1374 2513 1381 2516
rect 1374 2436 1377 2513
rect 1374 2433 1381 2436
rect 1378 2413 1381 2433
rect 1290 2326 1293 2346
rect 1298 2343 1301 2366
rect 1282 2323 1293 2326
rect 1282 2256 1285 2323
rect 1282 2253 1293 2256
rect 1178 2106 1181 2126
rect 1186 2113 1189 2126
rect 1194 2113 1197 2146
rect 1226 2143 1237 2146
rect 1234 2126 1237 2136
rect 1250 2126 1253 2216
rect 1266 2166 1269 2226
rect 1274 2213 1277 2226
rect 1274 2193 1277 2206
rect 1266 2163 1277 2166
rect 1210 2123 1221 2126
rect 1234 2123 1253 2126
rect 1210 2113 1221 2116
rect 1178 2103 1189 2106
rect 1226 2036 1229 2086
rect 1090 2033 1101 2036
rect 1218 2033 1229 2036
rect 1026 2013 1029 2026
rect 962 1983 989 1986
rect 890 1823 893 1836
rect 906 1823 917 1826
rect 906 1816 909 1823
rect 834 1793 837 1816
rect 874 1813 885 1816
rect 890 1813 909 1816
rect 714 1593 725 1596
rect 746 1593 749 1606
rect 754 1603 757 1616
rect 714 1533 717 1593
rect 722 1526 725 1586
rect 698 1433 701 1456
rect 666 1386 669 1406
rect 690 1393 693 1426
rect 706 1416 709 1526
rect 714 1523 725 1526
rect 738 1496 741 1546
rect 762 1533 765 1556
rect 762 1513 765 1526
rect 730 1493 741 1496
rect 714 1423 717 1446
rect 706 1413 725 1416
rect 730 1413 733 1493
rect 770 1446 773 1526
rect 762 1443 773 1446
rect 762 1416 765 1443
rect 770 1423 773 1436
rect 738 1406 741 1416
rect 762 1413 773 1416
rect 666 1383 685 1386
rect 610 1213 613 1266
rect 610 1103 613 1126
rect 578 1023 589 1026
rect 506 933 525 936
rect 498 913 501 926
rect 514 913 517 926
rect 530 906 533 926
rect 546 923 549 936
rect 470 883 485 886
rect 434 843 445 846
rect 434 813 437 836
rect 442 813 445 843
rect 426 736 429 796
rect 434 773 437 806
rect 466 803 469 816
rect 474 803 477 856
rect 426 733 453 736
rect 426 723 429 733
rect 466 723 469 796
rect 482 733 485 883
rect 506 846 509 906
rect 530 903 541 906
rect 506 843 517 846
rect 498 813 501 826
rect 514 813 517 843
rect 522 813 525 826
rect 546 823 549 916
rect 562 913 565 956
rect 570 913 573 936
rect 578 923 581 1016
rect 586 916 589 1023
rect 618 1013 621 1136
rect 626 1093 629 1136
rect 634 993 637 1176
rect 642 1113 645 1196
rect 650 1173 653 1346
rect 682 1266 685 1383
rect 682 1263 693 1266
rect 666 1213 669 1226
rect 690 1193 693 1263
rect 698 1233 701 1406
rect 730 1403 741 1406
rect 754 1403 765 1406
rect 706 1263 709 1336
rect 722 1333 725 1396
rect 714 1313 717 1326
rect 730 1323 733 1403
rect 738 1223 741 1336
rect 746 1296 749 1326
rect 754 1316 757 1386
rect 770 1333 773 1413
rect 754 1313 765 1316
rect 778 1303 781 1616
rect 786 1536 789 1726
rect 802 1723 805 1736
rect 810 1706 813 1736
rect 818 1723 821 1746
rect 842 1733 845 1746
rect 866 1736 869 1746
rect 806 1703 813 1706
rect 794 1543 797 1636
rect 806 1626 809 1703
rect 806 1623 813 1626
rect 786 1533 797 1536
rect 802 1533 805 1606
rect 810 1586 813 1623
rect 818 1603 821 1716
rect 834 1713 837 1726
rect 842 1713 845 1726
rect 850 1716 853 1736
rect 858 1733 869 1736
rect 858 1723 861 1733
rect 874 1726 877 1756
rect 866 1723 877 1726
rect 850 1713 861 1716
rect 826 1613 829 1626
rect 810 1583 817 1586
rect 786 1513 789 1526
rect 794 1496 797 1533
rect 790 1493 797 1496
rect 790 1426 793 1493
rect 790 1423 797 1426
rect 794 1406 797 1423
rect 786 1403 797 1406
rect 802 1393 805 1516
rect 814 1436 817 1583
rect 834 1546 837 1616
rect 826 1543 837 1546
rect 814 1433 821 1436
rect 810 1413 813 1426
rect 786 1323 797 1326
rect 786 1313 789 1323
rect 746 1293 753 1296
rect 750 1216 753 1293
rect 818 1243 821 1433
rect 826 1423 829 1543
rect 842 1523 845 1706
rect 858 1633 861 1713
rect 850 1556 853 1626
rect 866 1613 869 1626
rect 874 1623 877 1716
rect 882 1583 885 1736
rect 890 1606 893 1806
rect 898 1613 901 1636
rect 906 1623 909 1726
rect 914 1723 917 1816
rect 922 1753 925 1836
rect 930 1823 941 1826
rect 938 1813 941 1823
rect 930 1783 933 1806
rect 914 1703 917 1716
rect 930 1673 933 1736
rect 954 1726 957 1816
rect 962 1803 965 1946
rect 970 1933 973 1956
rect 970 1913 973 1926
rect 978 1803 981 1936
rect 986 1923 989 1983
rect 986 1813 989 1856
rect 994 1823 997 1936
rect 1010 1933 1013 1946
rect 1018 1903 1021 1916
rect 1026 1906 1029 1926
rect 1042 1923 1069 1926
rect 1026 1903 1033 1906
rect 1058 1903 1061 1916
rect 1010 1813 1013 1836
rect 1018 1813 1021 1886
rect 1030 1806 1033 1903
rect 1074 1833 1077 1936
rect 1082 1883 1085 2016
rect 1090 1986 1093 2033
rect 1106 2003 1109 2016
rect 1130 1993 1133 2016
rect 1090 1983 1109 1986
rect 1106 1933 1109 1983
rect 1162 1936 1165 1946
rect 1114 1926 1117 1936
rect 1146 1933 1165 1936
rect 1106 1916 1109 1926
rect 1114 1923 1141 1926
rect 1106 1913 1125 1916
rect 1122 1903 1125 1913
rect 1146 1903 1149 1933
rect 1154 1923 1165 1926
rect 1050 1813 1053 1826
rect 1114 1823 1117 1836
rect 1122 1833 1125 1886
rect 1154 1883 1157 1916
rect 1162 1876 1165 1923
rect 1170 1896 1173 1966
rect 1186 1943 1189 2016
rect 1194 1963 1197 2016
rect 1178 1923 1189 1926
rect 1178 1903 1181 1916
rect 1170 1893 1181 1896
rect 1178 1883 1181 1893
rect 1162 1873 1173 1876
rect 994 1793 997 1806
rect 1002 1803 1013 1806
rect 1026 1803 1033 1806
rect 954 1723 965 1726
rect 970 1723 973 1746
rect 1010 1733 1021 1736
rect 914 1613 917 1626
rect 890 1603 901 1606
rect 898 1573 901 1603
rect 850 1553 869 1556
rect 850 1533 853 1546
rect 834 1513 853 1516
rect 858 1446 861 1526
rect 866 1496 869 1553
rect 874 1513 877 1526
rect 866 1493 873 1496
rect 882 1493 885 1536
rect 890 1523 909 1526
rect 922 1523 925 1636
rect 930 1543 933 1626
rect 938 1566 941 1636
rect 954 1613 957 1646
rect 962 1633 965 1723
rect 938 1563 949 1566
rect 946 1523 949 1563
rect 970 1533 973 1626
rect 994 1603 997 1676
rect 1010 1643 1013 1733
rect 1018 1713 1021 1726
rect 1026 1723 1029 1803
rect 1098 1793 1101 1816
rect 1122 1813 1133 1816
rect 1138 1806 1141 1826
rect 1146 1813 1149 1866
rect 1162 1823 1165 1846
rect 1170 1816 1173 1873
rect 1194 1836 1197 1956
rect 1218 1946 1221 2033
rect 1218 1943 1229 1946
rect 1178 1833 1197 1836
rect 1162 1813 1173 1816
rect 1034 1696 1037 1736
rect 1026 1693 1037 1696
rect 1042 1693 1045 1726
rect 1026 1636 1029 1693
rect 1050 1673 1053 1736
rect 1066 1723 1069 1766
rect 1074 1733 1077 1746
rect 1082 1723 1085 1736
rect 1090 1703 1093 1736
rect 1106 1733 1117 1736
rect 1130 1733 1133 1806
rect 1138 1803 1149 1806
rect 1146 1743 1173 1746
rect 1106 1676 1109 1733
rect 1122 1683 1125 1726
rect 1082 1673 1109 1676
rect 1026 1633 1037 1636
rect 1034 1613 1037 1633
rect 986 1533 989 1546
rect 1034 1526 1037 1536
rect 954 1523 973 1526
rect 850 1443 861 1446
rect 842 1413 845 1426
rect 850 1333 853 1443
rect 858 1423 861 1436
rect 858 1333 861 1406
rect 870 1346 873 1493
rect 890 1466 893 1523
rect 882 1463 893 1466
rect 882 1413 885 1463
rect 930 1446 933 1516
rect 938 1503 941 1516
rect 954 1506 957 1523
rect 986 1516 989 1526
rect 962 1513 989 1516
rect 1010 1523 1037 1526
rect 1042 1523 1045 1646
rect 1074 1533 1077 1626
rect 1082 1603 1085 1673
rect 1090 1613 1093 1666
rect 1106 1613 1109 1636
rect 1138 1633 1141 1736
rect 1146 1733 1149 1743
rect 1146 1703 1149 1726
rect 1154 1723 1157 1736
rect 1170 1733 1173 1743
rect 1186 1736 1189 1826
rect 1202 1813 1205 1916
rect 1210 1863 1213 1916
rect 1218 1913 1221 1926
rect 1226 1906 1229 1943
rect 1234 1913 1237 2026
rect 1258 2016 1261 2136
rect 1274 2133 1277 2163
rect 1266 2073 1269 2106
rect 1274 2103 1277 2116
rect 1290 2113 1293 2253
rect 1298 2233 1301 2336
rect 1306 2283 1309 2336
rect 1314 2323 1317 2396
rect 1346 2393 1349 2406
rect 1386 2343 1389 2656
rect 1402 2616 1405 2763
rect 1394 2613 1405 2616
rect 1394 2393 1397 2613
rect 1402 2593 1405 2606
rect 1410 2526 1413 2616
rect 1402 2523 1413 2526
rect 1402 2513 1405 2523
rect 1418 2516 1421 2696
rect 1434 2623 1445 2626
rect 1426 2523 1429 2536
rect 1418 2513 1429 2516
rect 1434 2513 1437 2623
rect 1450 2613 1453 2726
rect 1482 2646 1485 2823
rect 1498 2813 1501 2866
rect 1490 2733 1493 2806
rect 1506 2756 1509 2836
rect 1498 2753 1509 2756
rect 1490 2713 1493 2726
rect 1498 2706 1501 2753
rect 1514 2746 1517 3040
rect 1530 3026 1533 3040
rect 1530 3023 1541 3026
rect 1538 2966 1541 3023
rect 1530 2963 1541 2966
rect 1530 2946 1533 2963
rect 1578 2946 1581 3040
rect 1594 3037 1613 3040
rect 1526 2943 1533 2946
rect 1526 2856 1529 2943
rect 1538 2933 1541 2946
rect 1578 2943 1605 2946
rect 1610 2943 1613 3037
rect 1850 3023 1853 3040
rect 1602 2936 1605 2943
rect 1526 2853 1533 2856
rect 1522 2823 1525 2836
rect 1474 2643 1485 2646
rect 1490 2703 1501 2706
rect 1506 2743 1517 2746
rect 1474 2603 1477 2643
rect 1490 2626 1493 2703
rect 1482 2623 1493 2626
rect 1490 2603 1493 2616
rect 1426 2413 1429 2513
rect 1442 2413 1445 2526
rect 1482 2523 1485 2536
rect 1490 2413 1493 2536
rect 1506 2523 1509 2743
rect 1514 2706 1517 2736
rect 1522 2723 1525 2816
rect 1530 2793 1533 2853
rect 1538 2833 1541 2916
rect 1562 2906 1565 2926
rect 1554 2903 1565 2906
rect 1554 2836 1557 2903
rect 1554 2833 1565 2836
rect 1562 2813 1565 2833
rect 1570 2813 1573 2926
rect 1578 2916 1581 2936
rect 1602 2933 1629 2936
rect 1626 2916 1629 2933
rect 1578 2913 1589 2916
rect 1586 2846 1589 2913
rect 1578 2843 1589 2846
rect 1618 2913 1629 2916
rect 1618 2846 1621 2913
rect 1618 2843 1629 2846
rect 1530 2733 1533 2766
rect 1538 2713 1541 2806
rect 1562 2796 1565 2806
rect 1546 2793 1565 2796
rect 1578 2763 1581 2843
rect 1586 2823 1621 2826
rect 1514 2703 1525 2706
rect 1522 2576 1525 2703
rect 1538 2583 1541 2616
rect 1546 2603 1549 2726
rect 1554 2643 1557 2736
rect 1570 2686 1573 2736
rect 1594 2723 1597 2806
rect 1610 2803 1613 2816
rect 1618 2766 1621 2823
rect 1626 2803 1629 2843
rect 1642 2826 1645 2936
rect 1682 2933 1685 2946
rect 1658 2916 1661 2926
rect 1666 2923 1677 2926
rect 1658 2913 1685 2916
rect 1690 2883 1693 2926
rect 1706 2906 1709 2926
rect 1722 2923 1725 2946
rect 1702 2903 1709 2906
rect 1702 2836 1705 2903
rect 1702 2833 1709 2836
rect 1634 2823 1645 2826
rect 1642 2803 1645 2823
rect 1658 2823 1685 2826
rect 1610 2763 1621 2766
rect 1610 2686 1613 2763
rect 1642 2693 1645 2776
rect 1650 2706 1653 2816
rect 1658 2813 1661 2823
rect 1666 2813 1685 2816
rect 1706 2813 1709 2833
rect 1658 2713 1661 2726
rect 1666 2716 1669 2806
rect 1674 2726 1677 2813
rect 1690 2803 1701 2806
rect 1706 2783 1709 2806
rect 1714 2773 1717 2886
rect 1722 2726 1725 2816
rect 1738 2803 1741 2916
rect 1770 2913 1773 2936
rect 1802 2856 1805 2956
rect 1882 2926 1885 3026
rect 1914 2956 1917 2976
rect 1922 2963 1925 3040
rect 2002 3037 2029 3040
rect 1906 2953 1925 2956
rect 1922 2933 1925 2953
rect 1802 2853 1809 2856
rect 1762 2803 1765 2816
rect 1674 2723 1709 2726
rect 1714 2723 1749 2726
rect 1666 2713 1677 2716
rect 1650 2703 1677 2706
rect 1570 2683 1589 2686
rect 1610 2683 1621 2686
rect 1570 2616 1573 2626
rect 1514 2573 1525 2576
rect 1514 2513 1517 2573
rect 1522 2413 1525 2526
rect 1538 2523 1541 2536
rect 1554 2503 1557 2616
rect 1562 2613 1573 2616
rect 1546 2426 1549 2436
rect 1538 2423 1549 2426
rect 1322 2313 1325 2326
rect 1298 2213 1301 2226
rect 1306 2223 1309 2236
rect 1298 2116 1301 2136
rect 1298 2113 1305 2116
rect 1250 2013 1261 2016
rect 1242 1993 1245 2006
rect 1226 1903 1237 1906
rect 1242 1893 1245 1916
rect 1250 1883 1253 2013
rect 1258 1993 1261 2006
rect 1282 2003 1285 2016
rect 1290 2013 1293 2076
rect 1302 2046 1305 2113
rect 1314 2103 1317 2296
rect 1322 2213 1325 2236
rect 1338 2213 1341 2226
rect 1346 2223 1349 2256
rect 1362 2213 1365 2226
rect 1370 2213 1373 2326
rect 1402 2236 1405 2376
rect 1418 2333 1421 2396
rect 1442 2393 1445 2406
rect 1426 2316 1429 2366
rect 1426 2313 1437 2316
rect 1386 2233 1405 2236
rect 1378 2213 1381 2226
rect 1346 2203 1365 2206
rect 1322 2133 1325 2156
rect 1330 2133 1333 2146
rect 1330 2123 1349 2126
rect 1330 2103 1333 2116
rect 1298 2043 1305 2046
rect 1298 2023 1301 2043
rect 1322 2013 1325 2026
rect 1346 2023 1349 2123
rect 1354 2063 1357 2156
rect 1362 2143 1365 2203
rect 1370 2193 1373 2206
rect 1386 2196 1389 2233
rect 1382 2193 1389 2196
rect 1370 2133 1373 2146
rect 1382 2136 1385 2193
rect 1394 2183 1397 2226
rect 1426 2213 1429 2306
rect 1402 2193 1405 2206
rect 1410 2173 1413 2206
rect 1434 2203 1437 2313
rect 1442 2303 1445 2326
rect 1378 2133 1385 2136
rect 1402 2133 1405 2156
rect 1378 2126 1381 2133
rect 1370 2123 1381 2126
rect 1258 1913 1261 1926
rect 1266 1913 1269 1966
rect 1202 1793 1205 1806
rect 1226 1803 1229 1816
rect 1178 1733 1189 1736
rect 1194 1733 1197 1776
rect 1226 1766 1229 1786
rect 1222 1763 1229 1766
rect 1178 1656 1181 1733
rect 1186 1723 1197 1726
rect 1202 1723 1205 1736
rect 1194 1706 1197 1723
rect 1194 1703 1201 1706
rect 954 1503 965 1506
rect 890 1423 893 1446
rect 922 1443 933 1446
rect 922 1413 925 1443
rect 930 1423 933 1436
rect 866 1343 873 1346
rect 866 1326 869 1343
rect 826 1306 829 1326
rect 850 1323 869 1326
rect 826 1303 845 1306
rect 746 1213 753 1216
rect 714 1193 717 1206
rect 650 1133 661 1136
rect 674 1133 677 1146
rect 658 1013 661 1116
rect 666 1023 669 1126
rect 674 1103 677 1126
rect 706 1076 709 1136
rect 722 1133 725 1176
rect 746 1143 749 1213
rect 762 1193 765 1216
rect 810 1196 813 1216
rect 802 1193 813 1196
rect 706 1073 717 1076
rect 714 1013 717 1073
rect 722 1013 725 1126
rect 746 1123 749 1136
rect 754 1116 757 1176
rect 802 1146 805 1193
rect 818 1173 821 1226
rect 826 1216 829 1296
rect 826 1213 845 1216
rect 834 1193 837 1206
rect 850 1203 853 1323
rect 882 1316 885 1396
rect 858 1313 885 1316
rect 858 1223 861 1306
rect 890 1246 893 1406
rect 898 1303 901 1336
rect 938 1333 941 1426
rect 946 1423 949 1446
rect 962 1403 965 1503
rect 1010 1456 1013 1523
rect 1034 1496 1037 1516
rect 1010 1453 1021 1456
rect 1002 1423 1005 1436
rect 970 1346 973 1406
rect 946 1343 973 1346
rect 922 1313 925 1326
rect 946 1323 949 1343
rect 962 1313 965 1326
rect 882 1243 893 1246
rect 858 1193 861 1206
rect 802 1143 813 1146
rect 746 1113 757 1116
rect 746 1026 749 1113
rect 802 1076 805 1126
rect 810 1086 813 1143
rect 818 1133 821 1146
rect 866 1133 869 1236
rect 874 1173 877 1216
rect 882 1213 885 1243
rect 970 1223 973 1336
rect 986 1333 989 1416
rect 994 1333 997 1406
rect 1010 1333 1013 1406
rect 1018 1326 1021 1453
rect 1026 1413 1029 1496
rect 1034 1493 1045 1496
rect 1042 1446 1045 1493
rect 1034 1443 1045 1446
rect 1034 1413 1037 1443
rect 1098 1413 1101 1606
rect 1122 1523 1125 1606
rect 1130 1603 1133 1616
rect 1138 1566 1141 1626
rect 1146 1586 1149 1656
rect 1170 1653 1181 1656
rect 1154 1593 1157 1606
rect 1146 1583 1157 1586
rect 1162 1583 1165 1606
rect 1154 1566 1157 1583
rect 1138 1563 1149 1566
rect 1154 1563 1161 1566
rect 1130 1533 1133 1556
rect 1130 1413 1133 1526
rect 1146 1523 1149 1563
rect 1158 1516 1161 1563
rect 1154 1513 1161 1516
rect 1138 1413 1141 1426
rect 1154 1406 1157 1513
rect 1170 1436 1173 1653
rect 1178 1613 1181 1646
rect 1186 1573 1189 1696
rect 1198 1616 1201 1703
rect 1194 1613 1201 1616
rect 1210 1613 1213 1736
rect 1222 1696 1225 1763
rect 1234 1703 1237 1746
rect 1222 1693 1229 1696
rect 1226 1616 1229 1693
rect 1242 1666 1245 1736
rect 1250 1683 1253 1816
rect 1266 1813 1269 1906
rect 1274 1903 1277 1926
rect 1306 1923 1309 2006
rect 1354 1923 1357 1936
rect 1370 1873 1373 2123
rect 1386 2113 1389 2126
rect 1402 2106 1405 2126
rect 1394 2103 1405 2106
rect 1386 2013 1389 2026
rect 1394 2003 1397 2103
rect 1426 2056 1429 2156
rect 1410 2053 1429 2056
rect 1386 1933 1389 1946
rect 1410 1943 1413 2053
rect 1434 2033 1437 2196
rect 1450 2156 1453 2246
rect 1458 2213 1461 2256
rect 1442 2153 1453 2156
rect 1466 2153 1469 2336
rect 1474 2203 1477 2226
rect 1482 2213 1485 2236
rect 1490 2213 1493 2326
rect 1498 2223 1501 2246
rect 1506 2223 1509 2236
rect 1530 2226 1533 2406
rect 1538 2333 1541 2423
rect 1554 2413 1557 2476
rect 1562 2413 1565 2613
rect 1570 2593 1573 2606
rect 1570 2533 1573 2546
rect 1570 2473 1573 2516
rect 1570 2423 1573 2446
rect 1514 2223 1533 2226
rect 1546 2223 1549 2406
rect 1570 2403 1573 2416
rect 1578 2413 1581 2506
rect 1586 2423 1589 2683
rect 1618 2626 1621 2683
rect 1618 2623 1629 2626
rect 1610 2593 1613 2616
rect 1626 2556 1629 2623
rect 1666 2613 1669 2646
rect 1674 2576 1677 2703
rect 1682 2693 1685 2706
rect 1698 2693 1701 2716
rect 1706 2713 1709 2723
rect 1714 2673 1717 2716
rect 1730 2623 1733 2716
rect 1738 2673 1741 2716
rect 1746 2713 1749 2723
rect 1754 2706 1757 2786
rect 1806 2766 1809 2853
rect 1818 2783 1821 2816
rect 1826 2803 1829 2926
rect 1866 2923 1885 2926
rect 1834 2823 1861 2826
rect 1802 2763 1809 2766
rect 1762 2713 1765 2726
rect 1770 2713 1773 2736
rect 1802 2733 1805 2763
rect 1850 2746 1853 2816
rect 1858 2813 1861 2823
rect 1858 2793 1861 2806
rect 1866 2803 1869 2923
rect 1882 2823 1885 2836
rect 1882 2793 1885 2806
rect 1834 2733 1837 2746
rect 1850 2743 1869 2746
rect 1778 2713 1781 2726
rect 1754 2703 1773 2706
rect 1682 2593 1685 2606
rect 1674 2573 1693 2576
rect 1618 2553 1629 2556
rect 1610 2523 1613 2546
rect 1618 2533 1621 2553
rect 1658 2523 1669 2526
rect 1666 2493 1669 2523
rect 1554 2326 1557 2336
rect 1562 2333 1565 2386
rect 1594 2376 1597 2446
rect 1626 2423 1629 2436
rect 1602 2393 1605 2406
rect 1578 2373 1597 2376
rect 1554 2323 1565 2326
rect 1578 2323 1581 2373
rect 1586 2306 1589 2366
rect 1610 2363 1613 2406
rect 1642 2403 1645 2426
rect 1666 2393 1669 2416
rect 1674 2413 1677 2526
rect 1682 2513 1685 2536
rect 1690 2533 1693 2573
rect 1698 2563 1701 2616
rect 1722 2596 1725 2616
rect 1714 2593 1725 2596
rect 1714 2533 1717 2593
rect 1690 2503 1693 2526
rect 1698 2523 1717 2526
rect 1722 2523 1725 2586
rect 1770 2583 1773 2646
rect 1778 2603 1781 2676
rect 1786 2613 1789 2626
rect 1786 2573 1789 2606
rect 1794 2593 1797 2716
rect 1818 2643 1821 2726
rect 1866 2696 1869 2743
rect 1882 2723 1885 2736
rect 1858 2693 1869 2696
rect 1858 2646 1861 2693
rect 1802 2576 1805 2636
rect 1810 2613 1813 2626
rect 1798 2573 1805 2576
rect 1746 2533 1749 2546
rect 1714 2423 1717 2516
rect 1578 2303 1589 2306
rect 1562 2223 1565 2246
rect 1578 2226 1581 2303
rect 1578 2223 1589 2226
rect 1442 2106 1445 2153
rect 1450 2123 1453 2146
rect 1482 2123 1485 2206
rect 1490 2133 1493 2146
rect 1498 2126 1501 2216
rect 1506 2203 1509 2216
rect 1514 2193 1517 2223
rect 1514 2133 1517 2166
rect 1490 2123 1501 2126
rect 1490 2113 1493 2123
rect 1442 2103 1449 2106
rect 1446 2016 1449 2103
rect 1442 2013 1449 2016
rect 1442 1993 1445 2013
rect 1458 1993 1461 2016
rect 1434 1913 1437 1926
rect 1474 1906 1477 1926
rect 1466 1903 1477 1906
rect 1258 1713 1261 1746
rect 1242 1663 1261 1666
rect 1222 1613 1229 1616
rect 1194 1593 1197 1613
rect 1222 1556 1225 1613
rect 1194 1533 1197 1546
rect 1210 1533 1213 1556
rect 1222 1553 1229 1556
rect 1226 1533 1229 1553
rect 1202 1513 1213 1516
rect 1218 1496 1221 1526
rect 1226 1506 1229 1526
rect 1234 1513 1237 1606
rect 1242 1563 1245 1616
rect 1250 1583 1253 1606
rect 1258 1603 1261 1663
rect 1266 1583 1269 1756
rect 1274 1693 1277 1766
rect 1282 1743 1285 1816
rect 1298 1813 1301 1826
rect 1306 1823 1317 1826
rect 1290 1763 1293 1806
rect 1306 1756 1309 1816
rect 1314 1773 1317 1823
rect 1290 1753 1309 1756
rect 1282 1723 1285 1736
rect 1290 1636 1293 1753
rect 1298 1736 1301 1746
rect 1298 1733 1309 1736
rect 1298 1713 1301 1726
rect 1306 1723 1309 1733
rect 1282 1633 1293 1636
rect 1282 1626 1285 1633
rect 1274 1623 1285 1626
rect 1290 1623 1301 1626
rect 1306 1623 1309 1706
rect 1274 1576 1277 1623
rect 1314 1616 1317 1736
rect 1322 1733 1325 1756
rect 1330 1736 1333 1826
rect 1338 1813 1349 1816
rect 1338 1783 1341 1813
rect 1330 1733 1341 1736
rect 1322 1703 1325 1726
rect 1330 1716 1333 1726
rect 1338 1723 1341 1733
rect 1346 1726 1349 1806
rect 1354 1803 1357 1816
rect 1362 1793 1365 1836
rect 1370 1813 1373 1866
rect 1394 1813 1397 1886
rect 1426 1813 1429 1836
rect 1434 1813 1437 1826
rect 1346 1723 1365 1726
rect 1330 1713 1341 1716
rect 1322 1623 1325 1646
rect 1330 1623 1333 1636
rect 1226 1503 1237 1506
rect 1218 1493 1229 1496
rect 1170 1433 1177 1436
rect 1034 1353 1037 1406
rect 1050 1363 1053 1406
rect 1138 1403 1157 1406
rect 1090 1346 1093 1366
rect 1026 1333 1029 1346
rect 898 1183 901 1206
rect 922 1193 925 1216
rect 810 1083 821 1086
rect 794 1073 805 1076
rect 794 1026 797 1073
rect 730 1023 749 1026
rect 730 1013 733 1023
rect 738 1006 741 1016
rect 722 956 725 1006
rect 690 953 725 956
rect 730 1003 741 1006
rect 602 933 613 936
rect 578 913 589 916
rect 594 923 605 926
rect 610 923 613 933
rect 626 923 629 936
rect 594 913 597 923
rect 554 806 557 906
rect 578 826 581 913
rect 586 836 589 906
rect 626 866 629 916
rect 610 863 629 866
rect 586 833 597 836
rect 562 813 565 826
rect 578 823 589 826
rect 570 813 581 816
rect 586 813 589 823
rect 514 733 517 806
rect 554 803 565 806
rect 530 726 533 736
rect 554 726 557 736
rect 514 723 533 726
rect 538 723 557 726
rect 562 716 565 796
rect 570 773 573 806
rect 586 733 589 806
rect 594 783 597 833
rect 594 723 597 736
rect 602 716 605 836
rect 610 823 613 863
rect 610 773 613 816
rect 618 813 621 856
rect 626 793 629 836
rect 634 823 637 936
rect 642 906 645 946
rect 658 923 661 936
rect 642 903 653 906
rect 658 883 661 916
rect 674 903 677 916
rect 682 883 685 916
rect 666 813 669 826
rect 682 823 685 836
rect 642 783 645 806
rect 690 796 693 953
rect 698 933 701 946
rect 698 913 701 926
rect 706 893 709 936
rect 722 933 725 946
rect 714 903 717 926
rect 730 923 733 1003
rect 746 996 749 1023
rect 762 1013 765 1026
rect 794 1023 805 1026
rect 738 993 749 996
rect 762 993 765 1006
rect 802 1003 805 1023
rect 722 856 725 876
rect 738 873 741 993
rect 810 983 813 1016
rect 818 1003 821 1083
rect 826 1013 829 1126
rect 842 1013 845 1036
rect 850 1013 853 1126
rect 866 1036 869 1126
rect 874 1103 877 1136
rect 906 1133 909 1176
rect 946 1133 949 1166
rect 898 1043 901 1126
rect 914 1113 917 1126
rect 866 1033 885 1036
rect 866 1013 869 1033
rect 874 1006 877 1026
rect 882 1016 885 1033
rect 890 1023 893 1036
rect 882 1013 893 1016
rect 842 1003 853 1006
rect 858 993 861 1006
rect 874 1003 885 1006
rect 746 933 749 956
rect 754 913 757 926
rect 698 803 701 816
rect 706 813 709 856
rect 718 853 725 856
rect 762 856 765 936
rect 778 933 781 966
rect 762 853 773 856
rect 706 796 709 806
rect 690 793 709 796
rect 442 703 445 716
rect 530 693 533 716
rect 546 713 565 716
rect 594 713 613 716
rect 618 713 621 726
rect 346 613 349 636
rect 418 626 421 636
rect 298 543 301 556
rect 306 533 309 546
rect 314 503 317 536
rect 322 523 325 606
rect 274 413 277 426
rect 210 323 221 326
rect 258 323 261 406
rect 282 403 285 436
rect 282 333 285 356
rect 290 333 293 416
rect 298 393 301 416
rect 322 403 325 416
rect 330 403 333 606
rect 338 603 349 606
rect 338 413 341 426
rect 346 406 349 603
rect 362 556 365 576
rect 358 553 365 556
rect 358 486 361 553
rect 370 496 373 546
rect 378 536 381 626
rect 394 613 397 626
rect 410 623 421 626
rect 434 623 445 626
rect 410 616 413 623
rect 402 613 413 616
rect 418 613 437 616
rect 402 593 405 606
rect 418 536 421 606
rect 442 556 445 623
rect 450 583 453 626
rect 466 623 477 626
rect 458 603 461 616
rect 466 573 469 623
rect 474 603 477 616
rect 434 553 445 556
rect 378 533 389 536
rect 418 533 429 536
rect 386 513 389 533
rect 394 523 405 526
rect 370 493 381 496
rect 358 483 365 486
rect 338 403 349 406
rect 314 383 317 396
rect 154 303 181 306
rect 130 193 133 216
rect 162 213 165 226
rect 170 183 173 206
rect 178 203 181 303
rect 202 213 205 236
rect 82 173 93 176
rect 90 133 93 173
rect 138 123 141 146
rect 186 143 189 206
rect 186 113 189 126
rect 202 123 205 206
rect 210 183 213 216
rect 218 213 221 323
rect 298 286 301 336
rect 314 326 317 336
rect 306 323 317 326
rect 322 323 325 376
rect 330 333 333 346
rect 314 306 317 323
rect 314 303 321 306
rect 298 283 309 286
rect 234 213 237 236
rect 226 193 229 206
rect 242 186 245 216
rect 258 203 261 226
rect 242 183 253 186
rect 250 143 253 183
rect 266 173 269 196
rect 282 193 285 226
rect 290 203 293 246
rect 298 203 301 256
rect 306 233 309 283
rect 318 236 321 303
rect 314 233 321 236
rect 258 133 261 146
rect 274 113 277 166
rect 298 156 301 176
rect 306 163 309 216
rect 314 203 317 233
rect 330 213 333 326
rect 338 236 341 403
rect 346 323 349 336
rect 338 233 349 236
rect 346 213 349 233
rect 298 153 309 156
rect 290 123 293 136
rect 306 133 309 153
rect 338 123 341 206
rect 362 173 365 483
rect 378 423 381 493
rect 386 486 389 506
rect 386 483 397 486
rect 394 426 397 483
rect 386 423 397 426
rect 378 393 381 416
rect 386 383 389 423
rect 402 393 405 406
rect 410 353 413 516
rect 418 513 421 526
rect 426 506 429 533
rect 434 523 437 553
rect 442 533 445 546
rect 426 503 437 506
rect 434 456 437 503
rect 426 453 437 456
rect 426 433 429 453
rect 426 413 429 426
rect 386 323 389 346
rect 450 343 453 406
rect 458 336 461 436
rect 466 403 469 536
rect 482 533 485 656
rect 490 603 493 626
rect 570 623 573 636
rect 618 633 621 706
rect 626 693 629 776
rect 666 733 669 746
rect 706 743 709 793
rect 718 786 721 853
rect 730 813 733 826
rect 770 813 773 853
rect 778 823 781 926
rect 718 783 725 786
rect 730 783 733 806
rect 722 763 725 783
rect 746 773 749 806
rect 722 733 725 756
rect 634 723 661 726
rect 634 653 637 723
rect 658 633 661 716
rect 642 623 661 626
rect 482 433 485 516
rect 490 503 493 526
rect 498 426 501 616
rect 522 593 525 606
rect 554 603 565 606
rect 562 536 565 603
rect 570 593 573 616
rect 586 573 589 606
rect 562 533 573 536
rect 506 513 509 526
rect 514 496 517 526
rect 522 506 525 526
rect 530 523 541 526
rect 538 513 557 516
rect 562 513 565 526
rect 522 503 533 506
rect 514 493 525 496
rect 482 423 501 426
rect 458 333 469 336
rect 386 113 389 206
rect 402 193 405 226
rect 410 213 429 216
rect 434 213 437 326
rect 442 296 445 326
rect 450 313 453 326
rect 466 316 469 333
rect 474 323 477 386
rect 482 333 485 423
rect 490 413 501 416
rect 506 413 509 436
rect 506 376 509 406
rect 498 373 509 376
rect 498 333 501 373
rect 514 336 517 426
rect 522 413 525 493
rect 530 393 533 436
rect 538 383 541 426
rect 546 423 549 436
rect 554 413 557 513
rect 570 493 573 533
rect 578 523 581 536
rect 586 513 589 536
rect 594 523 597 606
rect 626 603 637 606
rect 618 533 621 566
rect 602 506 605 526
rect 514 333 541 336
rect 514 323 517 333
rect 466 313 485 316
rect 498 303 501 316
rect 514 303 517 316
rect 538 313 541 326
rect 546 303 549 326
rect 562 323 565 436
rect 570 413 573 426
rect 578 423 581 506
rect 602 503 613 506
rect 586 413 589 436
rect 594 433 597 496
rect 610 446 613 503
rect 602 443 613 446
rect 602 423 605 443
rect 626 423 629 536
rect 634 513 637 526
rect 610 403 613 416
rect 570 323 573 336
rect 602 323 605 346
rect 642 343 645 606
rect 650 523 653 623
rect 658 613 661 623
rect 666 613 669 626
rect 658 593 661 606
rect 674 536 677 616
rect 682 606 685 636
rect 690 613 693 626
rect 698 613 701 716
rect 730 703 733 736
rect 746 733 749 746
rect 762 733 765 766
rect 738 713 741 726
rect 762 713 765 726
rect 682 603 701 606
rect 658 423 661 536
rect 674 533 685 536
rect 682 516 685 533
rect 674 513 685 516
rect 698 513 701 546
rect 666 443 669 506
rect 666 406 669 416
rect 674 413 677 513
rect 682 406 685 506
rect 690 423 693 496
rect 698 413 701 446
rect 706 433 709 616
rect 722 613 725 626
rect 714 583 717 606
rect 730 593 733 606
rect 746 603 749 696
rect 778 686 781 776
rect 794 773 797 936
rect 818 923 821 936
rect 826 806 829 926
rect 874 923 877 996
rect 882 976 885 1003
rect 890 993 893 1006
rect 882 973 893 976
rect 834 813 837 826
rect 826 803 845 806
rect 850 803 853 826
rect 874 793 877 806
rect 882 786 885 936
rect 890 923 893 973
rect 898 926 901 1006
rect 906 1003 909 1096
rect 906 933 909 976
rect 914 953 917 1016
rect 922 1003 925 1056
rect 930 1013 933 1116
rect 970 1076 973 1166
rect 962 1073 973 1076
rect 938 1013 941 1026
rect 898 923 909 926
rect 914 923 917 936
rect 922 923 925 936
rect 906 913 909 923
rect 930 916 933 1006
rect 962 976 965 1073
rect 978 1053 981 1326
rect 1010 1293 1013 1326
rect 1018 1323 1029 1326
rect 1026 1313 1029 1323
rect 1042 1306 1045 1336
rect 1066 1323 1069 1346
rect 1086 1343 1093 1346
rect 1018 1303 1045 1306
rect 1018 1286 1021 1303
rect 1010 1283 1021 1286
rect 978 1023 981 1046
rect 986 1013 989 1246
rect 994 1173 997 1216
rect 1010 1143 1013 1283
rect 1034 1213 1037 1226
rect 1042 1146 1045 1296
rect 1074 1183 1077 1336
rect 1086 1286 1089 1343
rect 1086 1283 1093 1286
rect 1090 1236 1093 1283
rect 1090 1233 1097 1236
rect 1082 1176 1085 1226
rect 1094 1186 1097 1233
rect 1106 1213 1109 1236
rect 1114 1213 1117 1296
rect 1122 1203 1125 1326
rect 1130 1306 1133 1336
rect 1146 1323 1149 1403
rect 1162 1386 1165 1426
rect 1174 1386 1177 1433
rect 1158 1383 1165 1386
rect 1170 1383 1177 1386
rect 1158 1326 1161 1383
rect 1170 1363 1173 1383
rect 1170 1333 1173 1356
rect 1158 1323 1165 1326
rect 1130 1303 1141 1306
rect 1138 1246 1141 1303
rect 1130 1243 1141 1246
rect 1130 1223 1133 1243
rect 1162 1233 1165 1323
rect 1186 1316 1189 1456
rect 1202 1413 1205 1426
rect 1194 1403 1205 1406
rect 1194 1323 1197 1396
rect 1202 1373 1205 1403
rect 1218 1386 1221 1416
rect 1226 1393 1229 1493
rect 1234 1413 1237 1503
rect 1218 1383 1229 1386
rect 1186 1313 1197 1316
rect 1130 1206 1133 1216
rect 1154 1213 1157 1226
rect 1130 1203 1141 1206
rect 1074 1173 1085 1176
rect 1090 1183 1097 1186
rect 1130 1183 1133 1196
rect 994 1113 997 1126
rect 978 993 981 1006
rect 986 983 989 1006
rect 1002 983 1005 1006
rect 1018 1003 1021 1076
rect 962 973 973 976
rect 938 923 941 936
rect 922 913 933 916
rect 946 913 949 956
rect 954 933 965 936
rect 922 896 925 913
rect 954 903 957 916
rect 914 893 925 896
rect 914 836 917 893
rect 938 856 941 896
rect 970 893 973 973
rect 978 933 981 966
rect 978 913 981 926
rect 934 853 941 856
rect 914 833 925 836
rect 922 813 925 833
rect 898 786 901 806
rect 874 783 885 786
rect 890 783 901 786
rect 802 723 805 746
rect 874 736 877 783
rect 882 743 885 756
rect 858 733 877 736
rect 858 723 861 733
rect 866 713 869 726
rect 882 713 885 726
rect 890 723 893 783
rect 898 726 901 776
rect 934 766 937 853
rect 978 846 981 906
rect 994 886 997 936
rect 1018 923 1021 936
rect 1026 903 1029 1146
rect 1034 1143 1045 1146
rect 1050 1143 1053 1156
rect 1034 1116 1037 1143
rect 1042 1133 1069 1136
rect 1042 1123 1045 1133
rect 1034 1113 1041 1116
rect 1050 1113 1053 1126
rect 1066 1123 1069 1133
rect 1038 1056 1041 1113
rect 1038 1053 1045 1056
rect 1034 1013 1037 1036
rect 1042 1003 1045 1053
rect 1050 1013 1053 1066
rect 1058 943 1061 1026
rect 1074 1016 1077 1173
rect 1090 1163 1093 1183
rect 1090 1133 1093 1146
rect 1082 1026 1085 1046
rect 1082 1023 1089 1026
rect 1098 1023 1101 1036
rect 1066 1013 1077 1016
rect 1066 936 1069 1013
rect 1058 933 1069 936
rect 1058 886 1061 933
rect 1074 923 1077 1006
rect 1086 946 1089 1023
rect 1098 963 1101 1016
rect 1106 953 1109 1006
rect 1114 1003 1117 1126
rect 1138 1123 1141 1203
rect 1154 1166 1157 1206
rect 1154 1163 1161 1166
rect 1170 1163 1173 1206
rect 1158 1086 1161 1163
rect 1154 1083 1161 1086
rect 1082 943 1089 946
rect 994 883 1005 886
rect 970 843 981 846
rect 954 793 957 816
rect 970 796 973 843
rect 1002 803 1005 883
rect 1050 883 1061 886
rect 1026 813 1029 826
rect 970 793 981 796
rect 934 763 941 766
rect 906 733 917 736
rect 922 733 925 746
rect 898 723 909 726
rect 914 723 917 733
rect 778 683 789 686
rect 770 613 773 626
rect 770 566 773 606
rect 786 576 789 683
rect 810 593 813 616
rect 858 613 869 616
rect 874 613 877 626
rect 890 603 893 626
rect 898 603 901 616
rect 922 606 925 726
rect 938 686 941 763
rect 962 713 965 726
rect 938 683 949 686
rect 930 613 933 626
rect 906 603 917 606
rect 922 603 933 606
rect 930 583 933 603
rect 786 573 805 576
rect 770 563 789 566
rect 746 533 749 556
rect 754 533 757 546
rect 770 533 773 546
rect 786 526 789 563
rect 802 556 805 573
rect 802 553 809 556
rect 746 523 765 526
rect 786 523 797 526
rect 722 493 725 516
rect 714 423 717 436
rect 738 423 749 426
rect 714 413 725 416
rect 666 403 685 406
rect 714 346 717 413
rect 722 356 725 406
rect 738 373 741 423
rect 754 416 757 446
rect 746 413 757 416
rect 762 413 765 436
rect 746 403 749 413
rect 754 383 757 406
rect 770 393 773 406
rect 722 353 733 356
rect 674 343 685 346
rect 714 343 725 346
rect 618 333 645 336
rect 442 293 453 296
rect 450 226 453 293
rect 442 223 453 226
rect 418 193 421 206
rect 426 143 429 213
rect 442 123 445 223
rect 458 163 461 206
rect 450 123 453 136
rect 466 113 469 216
rect 506 213 509 226
rect 514 223 517 246
rect 474 123 477 206
rect 522 156 525 236
rect 530 223 541 226
rect 530 206 533 216
rect 554 213 557 226
rect 562 213 565 226
rect 586 213 589 306
rect 594 213 597 316
rect 530 203 557 206
rect 514 153 525 156
rect 482 143 501 146
rect 482 133 485 143
rect 490 103 493 136
rect 498 113 501 143
rect 514 126 517 153
rect 522 136 525 146
rect 522 133 533 136
rect 514 123 525 126
rect 530 123 533 133
rect 538 123 541 196
rect 546 133 549 146
rect 554 136 557 203
rect 586 173 589 206
rect 602 166 605 226
rect 610 173 613 226
rect 618 213 621 333
rect 634 313 637 326
rect 666 313 669 336
rect 674 323 677 336
rect 682 276 685 343
rect 690 323 701 326
rect 666 273 685 276
rect 626 213 629 256
rect 626 166 629 176
rect 554 133 565 136
rect 562 123 565 133
rect 570 113 573 166
rect 602 163 629 166
rect 602 116 605 163
rect 634 143 637 206
rect 650 163 653 226
rect 658 213 661 226
rect 666 206 669 273
rect 698 266 701 316
rect 706 303 709 326
rect 722 313 725 343
rect 730 313 733 353
rect 714 283 717 306
rect 738 303 741 316
rect 674 223 677 266
rect 690 263 701 266
rect 682 216 685 226
rect 690 223 693 263
rect 674 213 685 216
rect 666 203 685 206
rect 682 143 685 203
rect 690 193 693 206
rect 626 133 637 136
rect 698 133 701 236
rect 706 223 709 246
rect 714 226 717 266
rect 714 223 733 226
rect 722 193 725 216
rect 730 213 733 223
rect 746 213 749 326
rect 730 156 733 206
rect 730 153 741 156
rect 706 133 709 146
rect 602 113 613 116
rect 642 113 645 126
rect 650 123 661 126
rect 698 113 701 126
rect 738 113 741 153
rect 754 123 757 316
rect 762 223 765 316
rect 770 293 773 326
rect 778 303 781 416
rect 786 413 789 516
rect 794 503 797 523
rect 806 496 809 553
rect 818 533 829 536
rect 818 513 821 526
rect 834 523 837 536
rect 850 533 853 566
rect 946 563 949 683
rect 970 603 973 616
rect 874 523 877 546
rect 802 493 809 496
rect 786 383 789 406
rect 802 403 805 493
rect 826 393 829 416
rect 834 386 837 436
rect 826 383 837 386
rect 842 383 845 506
rect 882 413 885 526
rect 930 523 933 536
rect 946 456 949 546
rect 978 543 981 793
rect 1018 783 1021 796
rect 1050 773 1053 883
rect 1082 833 1085 943
rect 1090 913 1093 926
rect 1098 816 1101 936
rect 1106 923 1109 946
rect 1122 936 1125 1016
rect 1138 1013 1141 1046
rect 1154 1006 1157 1083
rect 1170 1046 1173 1126
rect 1194 1056 1197 1313
rect 1202 1173 1205 1366
rect 1210 1316 1213 1336
rect 1210 1313 1217 1316
rect 1214 1236 1217 1313
rect 1226 1303 1229 1383
rect 1210 1233 1217 1236
rect 1210 1186 1213 1233
rect 1218 1193 1221 1216
rect 1210 1183 1221 1186
rect 1250 1183 1253 1536
rect 1258 1533 1261 1576
rect 1266 1573 1277 1576
rect 1282 1613 1309 1616
rect 1314 1613 1333 1616
rect 1266 1503 1269 1573
rect 1274 1423 1277 1526
rect 1282 1413 1285 1613
rect 1290 1553 1293 1606
rect 1306 1546 1309 1556
rect 1290 1543 1309 1546
rect 1290 1513 1293 1543
rect 1330 1533 1333 1586
rect 1338 1526 1341 1713
rect 1346 1703 1349 1716
rect 1362 1703 1365 1723
rect 1362 1626 1365 1646
rect 1358 1623 1365 1626
rect 1346 1603 1349 1616
rect 1358 1556 1361 1623
rect 1358 1553 1365 1556
rect 1370 1553 1373 1776
rect 1394 1733 1405 1736
rect 1378 1713 1381 1726
rect 1378 1613 1381 1626
rect 1386 1623 1389 1716
rect 1386 1603 1389 1616
rect 1394 1596 1397 1616
rect 1402 1613 1405 1726
rect 1410 1723 1413 1736
rect 1418 1633 1421 1806
rect 1442 1673 1445 1876
rect 1466 1846 1469 1903
rect 1466 1843 1477 1846
rect 1450 1803 1453 1816
rect 1458 1803 1461 1826
rect 1466 1753 1469 1816
rect 1410 1613 1421 1616
rect 1386 1593 1397 1596
rect 1362 1533 1365 1553
rect 1386 1533 1389 1593
rect 1410 1546 1413 1613
rect 1418 1593 1421 1606
rect 1410 1543 1421 1546
rect 1426 1543 1429 1616
rect 1434 1603 1437 1626
rect 1442 1603 1445 1616
rect 1450 1596 1453 1726
rect 1474 1636 1477 1843
rect 1482 1813 1485 1826
rect 1482 1766 1485 1806
rect 1490 1803 1493 2016
rect 1498 2006 1501 2106
rect 1506 2013 1509 2126
rect 1522 2103 1525 2216
rect 1530 2163 1533 2206
rect 1586 2203 1589 2223
rect 1594 2203 1597 2316
rect 1618 2313 1621 2326
rect 1538 2133 1541 2156
rect 1610 2133 1613 2216
rect 1618 2193 1621 2206
rect 1634 2153 1637 2276
rect 1666 2273 1669 2336
rect 1682 2313 1685 2326
rect 1706 2323 1709 2416
rect 1722 2413 1725 2516
rect 1730 2423 1733 2446
rect 1738 2413 1741 2426
rect 1746 2413 1749 2516
rect 1746 2343 1749 2406
rect 1754 2403 1757 2456
rect 1762 2406 1765 2566
rect 1786 2523 1789 2546
rect 1798 2496 1801 2573
rect 1810 2503 1813 2606
rect 1818 2603 1821 2626
rect 1826 2603 1829 2616
rect 1826 2556 1829 2586
rect 1842 2566 1845 2646
rect 1858 2643 1869 2646
rect 1834 2563 1845 2566
rect 1826 2553 1837 2556
rect 1798 2493 1805 2496
rect 1770 2413 1797 2416
rect 1802 2413 1805 2493
rect 1810 2443 1821 2446
rect 1818 2426 1821 2443
rect 1810 2423 1821 2426
rect 1826 2423 1829 2436
rect 1834 2416 1837 2553
rect 1842 2523 1845 2536
rect 1850 2533 1853 2566
rect 1866 2563 1869 2643
rect 1874 2533 1877 2616
rect 1890 2543 1893 2686
rect 1898 2656 1901 2816
rect 1906 2726 1909 2756
rect 1914 2733 1917 2806
rect 1922 2753 1925 2926
rect 1970 2856 1973 2926
rect 2002 2906 2005 3037
rect 1998 2903 2005 2906
rect 1970 2853 1989 2856
rect 1938 2823 1941 2836
rect 1938 2793 1941 2806
rect 1930 2733 1933 2746
rect 1906 2723 1917 2726
rect 1898 2653 1909 2656
rect 1906 2606 1909 2653
rect 1946 2623 1949 2636
rect 1954 2616 1957 2726
rect 1906 2603 1917 2606
rect 1882 2533 1893 2536
rect 1898 2533 1901 2576
rect 1850 2503 1853 2526
rect 1866 2523 1877 2526
rect 1818 2413 1837 2416
rect 1842 2413 1845 2436
rect 1850 2423 1853 2446
rect 1866 2423 1869 2436
rect 1874 2413 1877 2516
rect 1762 2403 1781 2406
rect 1802 2356 1805 2406
rect 1802 2353 1813 2356
rect 1514 2016 1517 2026
rect 1514 2013 1525 2016
rect 1530 2013 1533 2026
rect 1498 2003 1509 2006
rect 1506 1926 1509 2003
rect 1514 1993 1517 2006
rect 1506 1923 1517 1926
rect 1522 1923 1525 2013
rect 1538 1926 1541 2006
rect 1538 1923 1545 1926
rect 1498 1813 1501 1836
rect 1506 1803 1509 1916
rect 1514 1813 1517 1923
rect 1530 1863 1533 1916
rect 1542 1836 1545 1923
rect 1538 1833 1545 1836
rect 1522 1813 1525 1826
rect 1538 1816 1541 1833
rect 1530 1813 1541 1816
rect 1554 1813 1557 2006
rect 1562 1953 1565 2016
rect 1578 1916 1581 2026
rect 1586 2006 1589 2126
rect 1634 2013 1637 2136
rect 1658 2133 1661 2216
rect 1714 2213 1717 2336
rect 1730 2313 1733 2336
rect 1802 2326 1805 2346
rect 1738 2223 1741 2246
rect 1666 2113 1669 2166
rect 1682 2046 1685 2126
rect 1682 2043 1689 2046
rect 1586 2003 1605 2006
rect 1594 1933 1597 1946
rect 1570 1913 1581 1916
rect 1530 1806 1533 1813
rect 1522 1803 1533 1806
rect 1546 1803 1557 1806
rect 1562 1803 1565 1816
rect 1514 1776 1517 1796
rect 1530 1793 1533 1803
rect 1514 1773 1521 1776
rect 1482 1763 1501 1766
rect 1498 1723 1501 1763
rect 1474 1633 1485 1636
rect 1442 1593 1453 1596
rect 1298 1523 1309 1526
rect 1314 1523 1341 1526
rect 1354 1523 1365 1526
rect 1298 1506 1301 1523
rect 1306 1513 1317 1516
rect 1322 1513 1325 1523
rect 1298 1503 1309 1506
rect 1298 1413 1301 1426
rect 1306 1423 1309 1503
rect 1314 1413 1317 1436
rect 1322 1433 1325 1506
rect 1266 1306 1269 1336
rect 1290 1316 1293 1326
rect 1274 1313 1293 1316
rect 1266 1303 1277 1306
rect 1298 1303 1301 1406
rect 1322 1313 1325 1426
rect 1330 1406 1333 1426
rect 1338 1423 1341 1516
rect 1362 1513 1381 1516
rect 1386 1513 1389 1526
rect 1330 1403 1341 1406
rect 1346 1403 1349 1416
rect 1354 1403 1357 1416
rect 1362 1413 1365 1513
rect 1370 1493 1373 1506
rect 1370 1423 1381 1426
rect 1370 1406 1373 1423
rect 1386 1416 1389 1426
rect 1362 1403 1373 1406
rect 1378 1413 1389 1416
rect 1338 1326 1341 1386
rect 1334 1323 1341 1326
rect 1266 1213 1269 1226
rect 1274 1213 1277 1303
rect 1334 1246 1337 1323
rect 1334 1243 1341 1246
rect 1282 1213 1285 1226
rect 1274 1203 1285 1206
rect 1218 1143 1221 1183
rect 1282 1166 1285 1186
rect 1274 1163 1285 1166
rect 1290 1163 1293 1236
rect 1330 1216 1333 1226
rect 1202 1096 1205 1136
rect 1218 1113 1221 1126
rect 1202 1093 1213 1096
rect 1138 1003 1157 1006
rect 1162 1043 1173 1046
rect 1186 1053 1197 1056
rect 1162 1003 1165 1043
rect 1186 1036 1189 1053
rect 1210 1046 1213 1093
rect 1234 1086 1237 1136
rect 1258 1113 1261 1126
rect 1274 1086 1277 1163
rect 1298 1146 1301 1216
rect 1314 1213 1333 1216
rect 1338 1206 1341 1243
rect 1306 1193 1309 1206
rect 1330 1203 1341 1206
rect 1346 1206 1349 1316
rect 1354 1213 1357 1316
rect 1362 1313 1365 1403
rect 1370 1323 1373 1396
rect 1378 1303 1381 1413
rect 1386 1326 1389 1406
rect 1394 1383 1397 1536
rect 1402 1476 1405 1496
rect 1402 1473 1409 1476
rect 1406 1366 1409 1473
rect 1418 1423 1421 1543
rect 1426 1493 1429 1526
rect 1434 1446 1437 1566
rect 1442 1506 1445 1593
rect 1458 1523 1461 1626
rect 1442 1503 1453 1506
rect 1466 1503 1469 1616
rect 1482 1546 1485 1633
rect 1474 1543 1485 1546
rect 1474 1523 1477 1543
rect 1506 1523 1509 1756
rect 1518 1616 1521 1773
rect 1518 1613 1525 1616
rect 1514 1583 1517 1606
rect 1426 1443 1437 1446
rect 1426 1406 1429 1443
rect 1450 1436 1453 1503
rect 1474 1466 1477 1516
rect 1402 1363 1409 1366
rect 1422 1403 1429 1406
rect 1386 1323 1397 1326
rect 1386 1246 1389 1316
rect 1378 1243 1389 1246
rect 1362 1233 1373 1236
rect 1346 1203 1357 1206
rect 1362 1203 1365 1226
rect 1298 1143 1305 1146
rect 1234 1083 1253 1086
rect 1274 1083 1285 1086
rect 1182 1033 1189 1036
rect 1202 1043 1213 1046
rect 1122 933 1133 936
rect 1138 933 1141 946
rect 1130 926 1133 933
rect 1122 913 1125 926
rect 1130 923 1141 926
rect 1138 913 1141 923
rect 1146 846 1149 966
rect 1154 893 1157 926
rect 1162 913 1165 926
rect 1138 843 1149 846
rect 1082 813 1101 816
rect 1114 813 1117 826
rect 1130 766 1133 836
rect 1138 776 1141 843
rect 1170 836 1173 1016
rect 1182 976 1185 1033
rect 1202 1023 1205 1043
rect 1182 973 1189 976
rect 1186 846 1189 973
rect 1202 936 1205 1016
rect 1198 933 1205 936
rect 1226 933 1229 1016
rect 1250 1003 1253 1083
rect 1266 956 1269 1026
rect 1282 996 1285 1083
rect 1302 1036 1305 1143
rect 1322 1133 1325 1166
rect 1302 1033 1309 1036
rect 1290 1003 1293 1026
rect 1282 993 1293 996
rect 1266 953 1277 956
rect 1198 876 1201 933
rect 1210 883 1213 926
rect 1258 906 1261 936
rect 1274 933 1277 953
rect 1290 913 1293 993
rect 1258 903 1269 906
rect 1198 873 1205 876
rect 1186 843 1193 846
rect 1170 833 1181 836
rect 1162 783 1165 816
rect 1178 776 1181 833
rect 1190 796 1193 843
rect 1138 773 1157 776
rect 1010 656 1013 726
rect 1018 723 1021 746
rect 1050 733 1053 766
rect 1130 763 1141 766
rect 1010 653 1017 656
rect 890 413 893 426
rect 898 396 901 416
rect 906 403 909 436
rect 914 403 917 456
rect 938 453 949 456
rect 898 393 917 396
rect 794 333 797 376
rect 802 313 805 346
rect 810 313 813 336
rect 818 303 821 326
rect 786 213 789 286
rect 826 283 829 383
rect 834 293 837 326
rect 802 223 813 226
rect 794 206 797 216
rect 762 103 765 206
rect 770 156 773 206
rect 786 203 797 206
rect 786 193 789 203
rect 802 193 805 223
rect 818 213 821 266
rect 842 236 845 316
rect 850 303 853 326
rect 858 303 861 316
rect 866 313 869 326
rect 826 233 845 236
rect 826 223 829 233
rect 834 163 837 226
rect 842 223 845 233
rect 858 226 861 286
rect 858 223 869 226
rect 770 153 781 156
rect 770 123 773 146
rect 778 133 781 153
rect 810 136 813 146
rect 794 133 805 136
rect 810 133 821 136
rect 826 133 829 146
rect 842 133 845 216
rect 858 203 861 223
rect 874 213 877 336
rect 898 326 901 336
rect 882 213 885 326
rect 890 323 901 326
rect 906 323 909 336
rect 914 323 917 393
rect 922 376 925 416
rect 938 403 941 453
rect 922 373 933 376
rect 922 333 925 366
rect 930 323 933 373
rect 890 303 893 323
rect 778 103 781 126
rect 810 113 813 126
rect 818 123 821 133
rect 866 106 869 206
rect 882 133 885 146
rect 882 113 885 126
rect 890 113 893 226
rect 898 223 901 316
rect 938 256 941 386
rect 946 333 949 346
rect 962 333 965 416
rect 970 363 973 526
rect 986 456 989 576
rect 1014 546 1017 653
rect 1026 593 1029 616
rect 1034 613 1037 626
rect 1042 613 1045 726
rect 1058 716 1061 726
rect 1066 723 1069 736
rect 1098 733 1109 736
rect 1138 733 1141 763
rect 1058 713 1077 716
rect 1042 593 1045 606
rect 1050 603 1053 616
rect 1058 576 1061 626
rect 1066 603 1069 616
rect 1010 543 1017 546
rect 1042 573 1061 576
rect 1010 513 1013 543
rect 1026 533 1037 536
rect 982 453 989 456
rect 982 406 985 453
rect 982 403 989 406
rect 978 333 981 386
rect 954 306 957 326
rect 986 316 989 403
rect 1018 396 1021 526
rect 1026 453 1029 526
rect 1026 403 1029 426
rect 1034 413 1037 526
rect 1042 523 1045 573
rect 1074 566 1077 713
rect 1090 706 1093 726
rect 1122 713 1125 726
rect 1090 703 1101 706
rect 1098 646 1101 703
rect 1130 686 1133 726
rect 1146 723 1149 746
rect 1154 736 1157 773
rect 1170 773 1181 776
rect 1186 793 1193 796
rect 1186 773 1189 793
rect 1154 733 1165 736
rect 1170 723 1173 773
rect 1194 733 1197 746
rect 1202 726 1205 873
rect 1194 723 1205 726
rect 1210 723 1213 826
rect 1242 823 1245 896
rect 1266 816 1269 903
rect 1298 886 1301 1016
rect 1306 1003 1309 1033
rect 1314 1023 1317 1126
rect 1330 1103 1333 1126
rect 1338 1023 1341 1136
rect 1354 1133 1357 1203
rect 1370 1196 1373 1233
rect 1378 1203 1381 1243
rect 1394 1236 1397 1323
rect 1386 1233 1397 1236
rect 1386 1223 1389 1233
rect 1402 1226 1405 1363
rect 1422 1346 1425 1403
rect 1410 1306 1413 1346
rect 1418 1343 1425 1346
rect 1418 1323 1421 1343
rect 1410 1303 1417 1306
rect 1434 1303 1437 1436
rect 1442 1433 1453 1436
rect 1466 1463 1477 1466
rect 1442 1403 1445 1433
rect 1450 1396 1453 1416
rect 1466 1406 1469 1463
rect 1482 1453 1485 1516
rect 1522 1483 1525 1613
rect 1530 1533 1533 1686
rect 1538 1603 1541 1626
rect 1546 1596 1549 1636
rect 1554 1623 1557 1803
rect 1562 1733 1565 1796
rect 1570 1763 1573 1826
rect 1578 1723 1581 1816
rect 1586 1716 1589 1826
rect 1594 1813 1597 1926
rect 1602 1883 1605 1926
rect 1602 1776 1605 1816
rect 1562 1703 1565 1716
rect 1578 1713 1589 1716
rect 1598 1773 1605 1776
rect 1562 1616 1565 1636
rect 1570 1623 1573 1646
rect 1578 1616 1581 1713
rect 1598 1706 1601 1773
rect 1594 1703 1601 1706
rect 1554 1613 1565 1616
rect 1570 1613 1581 1616
rect 1546 1593 1553 1596
rect 1538 1533 1541 1586
rect 1550 1516 1553 1593
rect 1562 1536 1565 1613
rect 1562 1533 1573 1536
rect 1546 1513 1553 1516
rect 1546 1493 1549 1513
rect 1562 1496 1565 1526
rect 1558 1493 1565 1496
rect 1558 1436 1561 1493
rect 1570 1446 1573 1533
rect 1578 1526 1581 1613
rect 1586 1536 1589 1626
rect 1594 1613 1597 1703
rect 1602 1603 1605 1616
rect 1610 1593 1613 1986
rect 1642 1956 1645 2006
rect 1658 1973 1661 2026
rect 1686 1996 1689 2043
rect 1682 1993 1689 1996
rect 1682 1976 1685 1993
rect 1698 1986 1701 2156
rect 1714 2133 1717 2156
rect 1722 2056 1725 2186
rect 1730 2163 1733 2216
rect 1730 2096 1733 2136
rect 1738 2123 1741 2136
rect 1746 2133 1749 2216
rect 1754 2126 1757 2216
rect 1762 2213 1765 2326
rect 1798 2323 1805 2326
rect 1762 2193 1765 2206
rect 1746 2123 1757 2126
rect 1746 2113 1749 2123
rect 1730 2093 1741 2096
rect 1722 2053 1729 2056
rect 1706 1993 1709 2016
rect 1698 1983 1709 1986
rect 1666 1973 1685 1976
rect 1642 1953 1653 1956
rect 1618 1903 1621 1936
rect 1626 1923 1629 1946
rect 1634 1813 1637 1936
rect 1650 1933 1653 1953
rect 1658 1923 1661 1936
rect 1666 1923 1669 1973
rect 1706 1966 1709 1983
rect 1726 1976 1729 2053
rect 1738 2013 1741 2093
rect 1762 2056 1765 2136
rect 1770 2133 1773 2186
rect 1778 2116 1781 2316
rect 1798 2256 1801 2323
rect 1798 2253 1805 2256
rect 1754 2053 1765 2056
rect 1774 2113 1781 2116
rect 1754 2013 1757 2053
rect 1774 2046 1777 2113
rect 1774 2043 1781 2046
rect 1778 2023 1781 2043
rect 1722 1973 1729 1976
rect 1706 1963 1713 1966
rect 1682 1846 1685 1936
rect 1710 1896 1713 1963
rect 1706 1893 1713 1896
rect 1722 1893 1725 1973
rect 1730 1923 1733 1946
rect 1746 1923 1749 2006
rect 1762 1993 1765 2006
rect 1770 1973 1773 2016
rect 1778 2003 1781 2016
rect 1786 2013 1789 2136
rect 1794 2133 1797 2156
rect 1762 1923 1765 1966
rect 1674 1843 1693 1846
rect 1674 1803 1677 1843
rect 1618 1733 1637 1736
rect 1626 1706 1629 1733
rect 1634 1713 1637 1726
rect 1642 1713 1645 1726
rect 1650 1716 1653 1766
rect 1658 1723 1661 1746
rect 1666 1733 1669 1766
rect 1650 1713 1661 1716
rect 1666 1713 1669 1726
rect 1690 1723 1693 1806
rect 1698 1743 1701 1816
rect 1626 1703 1637 1706
rect 1626 1603 1629 1616
rect 1634 1603 1637 1703
rect 1698 1646 1701 1716
rect 1706 1713 1709 1893
rect 1714 1816 1717 1866
rect 1714 1813 1733 1816
rect 1714 1783 1717 1806
rect 1722 1733 1725 1806
rect 1730 1713 1733 1813
rect 1738 1733 1741 1816
rect 1746 1813 1749 1826
rect 1754 1793 1757 1806
rect 1762 1776 1765 1836
rect 1770 1813 1773 1936
rect 1778 1923 1781 1996
rect 1786 1933 1789 2006
rect 1794 1993 1797 2126
rect 1802 2103 1805 2253
rect 1810 2193 1813 2353
rect 1818 2303 1821 2413
rect 1826 2256 1829 2346
rect 1842 2266 1845 2326
rect 1850 2316 1853 2406
rect 1866 2343 1869 2406
rect 1874 2393 1877 2406
rect 1858 2326 1861 2336
rect 1882 2333 1885 2466
rect 1890 2403 1893 2526
rect 1906 2523 1909 2596
rect 1914 2556 1917 2603
rect 1922 2593 1925 2616
rect 1930 2563 1933 2616
rect 1946 2613 1957 2616
rect 1962 2613 1965 2636
rect 1938 2593 1941 2606
rect 1946 2603 1949 2613
rect 1970 2603 1973 2816
rect 1986 2803 1989 2853
rect 1998 2826 2001 2903
rect 1998 2823 2005 2826
rect 2002 2803 2005 2823
rect 2010 2793 2013 2936
rect 2026 2933 2037 2936
rect 2050 2933 2053 2946
rect 2018 2823 2021 2836
rect 2026 2816 2029 2926
rect 2050 2903 2053 2916
rect 2066 2853 2069 2976
rect 2098 2956 2101 3040
rect 2146 2966 2149 3040
rect 2146 2963 2157 2966
rect 2098 2953 2109 2956
rect 2090 2923 2093 2946
rect 2106 2896 2109 2953
rect 2154 2933 2157 2963
rect 2162 2933 2173 2936
rect 2162 2903 2165 2926
rect 2170 2913 2181 2916
rect 2090 2893 2109 2896
rect 2058 2823 2061 2836
rect 2018 2813 2029 2816
rect 2010 2676 2013 2726
rect 2018 2723 2021 2813
rect 2026 2793 2029 2806
rect 2034 2753 2037 2816
rect 2090 2813 2093 2893
rect 2170 2866 2173 2913
rect 2170 2863 2181 2866
rect 2058 2793 2061 2806
rect 2122 2793 2125 2816
rect 2170 2803 2173 2856
rect 2178 2833 2181 2863
rect 2186 2766 2189 2926
rect 2194 2803 2197 2936
rect 2210 2933 2213 2946
rect 2226 2933 2229 2996
rect 2266 2966 2269 3040
rect 2282 2993 2285 3040
rect 2242 2963 2269 2966
rect 2418 2966 2421 3040
rect 2418 2963 2429 2966
rect 2202 2913 2213 2916
rect 2242 2886 2245 2963
rect 2266 2923 2269 2946
rect 2242 2883 2253 2886
rect 2234 2823 2237 2836
rect 2182 2763 2189 2766
rect 2026 2723 2029 2736
rect 2042 2733 2045 2746
rect 2002 2673 2013 2676
rect 1914 2553 1933 2556
rect 1914 2516 1917 2546
rect 1922 2523 1925 2536
rect 1914 2513 1925 2516
rect 1898 2403 1901 2446
rect 1930 2443 1933 2553
rect 1938 2533 1941 2546
rect 1946 2533 1949 2556
rect 1978 2546 1981 2626
rect 1986 2603 1989 2656
rect 1994 2603 1997 2616
rect 2002 2603 2005 2673
rect 2010 2596 2013 2656
rect 2018 2623 2029 2626
rect 2018 2603 2021 2616
rect 1994 2593 2013 2596
rect 1970 2543 1981 2546
rect 1954 2533 1965 2536
rect 1970 2526 1973 2543
rect 1978 2533 1981 2543
rect 1954 2503 1957 2526
rect 1962 2523 1973 2526
rect 1978 2483 1981 2526
rect 1986 2476 1989 2546
rect 1994 2503 1997 2593
rect 2026 2546 2029 2623
rect 2010 2543 2029 2546
rect 2002 2523 2005 2536
rect 1986 2473 1997 2476
rect 1914 2383 1917 2406
rect 1938 2393 1941 2416
rect 1994 2413 1997 2473
rect 2010 2413 2013 2543
rect 2034 2536 2037 2636
rect 2042 2613 2045 2726
rect 2058 2586 2061 2636
rect 2066 2613 2069 2726
rect 2074 2633 2077 2756
rect 2074 2613 2077 2626
rect 2074 2596 2077 2606
rect 2082 2603 2085 2676
rect 2090 2613 2093 2666
rect 2098 2606 2101 2626
rect 2106 2613 2109 2656
rect 2114 2606 2117 2636
rect 2122 2623 2125 2726
rect 2138 2686 2141 2746
rect 2138 2683 2149 2686
rect 2090 2603 2101 2606
rect 2106 2603 2117 2606
rect 2090 2596 2093 2603
rect 2106 2596 2109 2603
rect 2074 2593 2093 2596
rect 2098 2593 2109 2596
rect 2058 2583 2077 2586
rect 2018 2493 2021 2536
rect 2034 2533 2045 2536
rect 2050 2533 2069 2536
rect 2034 2506 2037 2526
rect 2042 2523 2045 2533
rect 2034 2503 2045 2506
rect 2050 2503 2053 2526
rect 2018 2423 2021 2436
rect 2034 2416 2037 2496
rect 2042 2463 2045 2503
rect 2066 2476 2069 2533
rect 2074 2493 2077 2583
rect 2082 2486 2085 2536
rect 2098 2523 2101 2593
rect 2114 2586 2117 2596
rect 2122 2593 2125 2606
rect 2106 2583 2117 2586
rect 2106 2523 2109 2583
rect 2138 2543 2141 2616
rect 2146 2563 2149 2683
rect 2154 2613 2157 2656
rect 2162 2623 2165 2636
rect 2170 2616 2173 2726
rect 2182 2686 2185 2763
rect 2182 2683 2189 2686
rect 2162 2613 2173 2616
rect 2154 2593 2157 2606
rect 2162 2603 2165 2613
rect 2178 2583 2181 2616
rect 2186 2613 2189 2683
rect 2202 2613 2205 2696
rect 2202 2593 2205 2606
rect 2082 2483 2093 2486
rect 2066 2473 2085 2476
rect 2042 2423 2045 2456
rect 2050 2423 2077 2426
rect 2034 2413 2045 2416
rect 2050 2413 2053 2423
rect 1858 2323 1885 2326
rect 1850 2313 1861 2316
rect 1858 2296 1861 2313
rect 1858 2293 1869 2296
rect 1842 2263 1853 2266
rect 1826 2253 1845 2256
rect 1810 2056 1813 2146
rect 1818 2133 1821 2216
rect 1826 2133 1829 2176
rect 1842 2126 1845 2253
rect 1850 2153 1853 2263
rect 1866 2236 1869 2293
rect 1858 2233 1869 2236
rect 1858 2173 1861 2233
rect 1866 2203 1869 2216
rect 1882 2213 1885 2323
rect 1898 2286 1901 2336
rect 1898 2283 1909 2286
rect 1858 2133 1861 2166
rect 1826 2123 1845 2126
rect 1826 2106 1829 2123
rect 1802 2053 1813 2056
rect 1822 2103 1829 2106
rect 1834 2113 1845 2116
rect 1802 1976 1805 2053
rect 1822 2036 1825 2103
rect 1822 2033 1829 2036
rect 1818 2003 1821 2016
rect 1794 1913 1797 1976
rect 1802 1973 1813 1976
rect 1810 1936 1813 1973
rect 1802 1903 1805 1936
rect 1810 1933 1821 1936
rect 1754 1773 1765 1776
rect 1770 1773 1773 1806
rect 1746 1733 1749 1756
rect 1754 1723 1757 1773
rect 1762 1706 1765 1736
rect 1770 1723 1773 1736
rect 1650 1633 1653 1646
rect 1690 1643 1701 1646
rect 1754 1703 1765 1706
rect 1618 1583 1621 1596
rect 1586 1533 1597 1536
rect 1602 1533 1605 1546
rect 1594 1526 1597 1533
rect 1578 1523 1589 1526
rect 1594 1523 1605 1526
rect 1586 1513 1589 1523
rect 1602 1513 1605 1523
rect 1610 1513 1613 1526
rect 1618 1523 1621 1576
rect 1626 1563 1629 1596
rect 1570 1443 1577 1446
rect 1474 1423 1477 1436
rect 1558 1433 1565 1436
rect 1474 1413 1493 1416
rect 1466 1403 1477 1406
rect 1450 1393 1461 1396
rect 1498 1393 1501 1406
rect 1442 1313 1445 1326
rect 1458 1323 1461 1393
rect 1466 1323 1477 1326
rect 1482 1323 1485 1336
rect 1490 1333 1493 1346
rect 1414 1246 1417 1303
rect 1394 1223 1405 1226
rect 1410 1243 1417 1246
rect 1362 1193 1373 1196
rect 1386 1193 1389 1206
rect 1362 1133 1365 1193
rect 1346 1123 1365 1126
rect 1394 1113 1397 1223
rect 1402 1143 1405 1216
rect 1410 1213 1413 1243
rect 1402 1093 1405 1116
rect 1410 1056 1413 1106
rect 1402 1053 1413 1056
rect 1314 936 1317 1016
rect 1322 983 1325 1006
rect 1306 933 1317 936
rect 1322 933 1325 946
rect 1330 933 1333 1006
rect 1306 906 1309 933
rect 1338 926 1341 1016
rect 1362 1003 1365 1016
rect 1386 1013 1389 1026
rect 1314 913 1317 926
rect 1330 923 1341 926
rect 1306 903 1321 906
rect 1298 883 1309 886
rect 1218 813 1245 816
rect 1266 813 1277 816
rect 1290 813 1301 816
rect 1218 803 1221 813
rect 1218 733 1221 756
rect 1090 643 1101 646
rect 1122 683 1133 686
rect 1090 613 1093 643
rect 1122 613 1125 683
rect 1138 613 1157 616
rect 1082 573 1085 606
rect 1090 593 1093 606
rect 1050 533 1053 566
rect 1058 563 1077 566
rect 1042 403 1045 516
rect 1058 476 1061 563
rect 1066 523 1069 536
rect 1050 473 1061 476
rect 1050 413 1053 473
rect 1066 423 1069 446
rect 1010 393 1021 396
rect 1010 333 1013 393
rect 1026 333 1029 356
rect 1058 353 1061 406
rect 1066 393 1069 406
rect 1066 346 1069 366
rect 1034 333 1037 346
rect 1058 343 1069 346
rect 978 313 989 316
rect 994 323 1013 326
rect 954 303 965 306
rect 930 253 941 256
rect 906 213 909 226
rect 914 213 917 236
rect 930 196 933 253
rect 962 246 965 303
rect 946 203 949 246
rect 954 243 965 246
rect 954 216 957 243
rect 978 236 981 313
rect 978 233 989 236
rect 954 213 973 216
rect 930 193 941 196
rect 978 193 981 206
rect 906 133 909 166
rect 938 163 941 193
rect 938 133 941 146
rect 914 123 933 126
rect 954 123 957 166
rect 914 113 917 123
rect 986 113 989 233
rect 994 213 997 323
rect 1034 303 1037 316
rect 1058 313 1061 343
rect 1074 323 1077 546
rect 1082 513 1085 556
rect 1106 533 1109 606
rect 1114 593 1117 606
rect 1122 536 1125 586
rect 1130 543 1133 606
rect 1122 533 1133 536
rect 1154 533 1157 613
rect 1170 603 1173 616
rect 1082 403 1085 416
rect 1090 363 1093 426
rect 1130 423 1133 533
rect 1162 523 1165 536
rect 1178 533 1181 586
rect 1194 576 1197 723
rect 1234 716 1237 813
rect 1242 793 1245 806
rect 1250 753 1253 806
rect 1274 803 1277 813
rect 1306 803 1309 883
rect 1250 723 1253 736
rect 1234 713 1253 716
rect 1218 603 1221 636
rect 1234 603 1237 636
rect 1242 596 1245 706
rect 1258 666 1261 726
rect 1274 716 1277 786
rect 1282 733 1285 796
rect 1290 733 1293 756
rect 1318 746 1321 903
rect 1330 753 1333 923
rect 1346 916 1349 926
rect 1354 923 1357 936
rect 1362 916 1365 926
rect 1346 913 1365 916
rect 1346 836 1349 913
rect 1338 833 1349 836
rect 1338 793 1341 833
rect 1370 823 1373 936
rect 1386 933 1389 966
rect 1402 956 1405 1053
rect 1426 1013 1429 1286
rect 1450 1193 1453 1216
rect 1442 1133 1445 1176
rect 1450 1116 1453 1146
rect 1442 1113 1453 1116
rect 1442 956 1445 1113
rect 1458 1096 1461 1296
rect 1466 1286 1469 1323
rect 1474 1303 1477 1316
rect 1490 1313 1493 1326
rect 1466 1283 1473 1286
rect 1470 1146 1473 1283
rect 1498 1233 1501 1356
rect 1506 1293 1509 1416
rect 1514 1353 1517 1406
rect 1522 1386 1525 1416
rect 1554 1393 1557 1416
rect 1522 1383 1533 1386
rect 1514 1333 1517 1346
rect 1530 1333 1533 1383
rect 1514 1313 1517 1326
rect 1522 1293 1525 1326
rect 1546 1283 1549 1366
rect 1562 1353 1565 1433
rect 1574 1356 1577 1443
rect 1602 1363 1605 1506
rect 1634 1456 1637 1596
rect 1642 1563 1645 1616
rect 1650 1573 1653 1626
rect 1658 1613 1661 1626
rect 1658 1523 1661 1546
rect 1630 1453 1637 1456
rect 1618 1403 1621 1416
rect 1630 1376 1633 1453
rect 1666 1426 1669 1556
rect 1682 1523 1685 1626
rect 1690 1606 1693 1643
rect 1754 1636 1757 1703
rect 1698 1613 1701 1636
rect 1754 1633 1765 1636
rect 1762 1613 1765 1633
rect 1690 1603 1701 1606
rect 1690 1553 1693 1603
rect 1714 1556 1717 1606
rect 1706 1553 1717 1556
rect 1706 1533 1709 1553
rect 1722 1533 1725 1566
rect 1738 1533 1741 1606
rect 1762 1533 1765 1546
rect 1762 1513 1765 1526
rect 1770 1523 1773 1566
rect 1662 1423 1669 1426
rect 1626 1373 1633 1376
rect 1574 1353 1581 1356
rect 1570 1323 1573 1346
rect 1578 1316 1581 1353
rect 1570 1313 1581 1316
rect 1570 1296 1573 1313
rect 1562 1293 1573 1296
rect 1490 1213 1509 1216
rect 1466 1143 1473 1146
rect 1466 1123 1469 1143
rect 1474 1113 1477 1126
rect 1482 1123 1485 1146
rect 1490 1133 1493 1213
rect 1522 1183 1525 1206
rect 1530 1143 1533 1176
rect 1538 1133 1541 1156
rect 1454 1093 1461 1096
rect 1454 1006 1457 1093
rect 1466 1013 1469 1106
rect 1454 1003 1461 1006
rect 1402 953 1413 956
rect 1386 893 1389 926
rect 1394 923 1397 936
rect 1410 933 1413 953
rect 1418 933 1421 956
rect 1442 953 1453 956
rect 1450 933 1453 953
rect 1458 933 1461 1003
rect 1474 996 1477 1026
rect 1470 993 1477 996
rect 1470 936 1473 993
rect 1470 933 1477 936
rect 1346 793 1349 816
rect 1386 806 1389 816
rect 1394 813 1397 886
rect 1402 846 1405 926
rect 1418 903 1421 926
rect 1426 893 1429 926
rect 1442 846 1445 926
rect 1458 903 1461 926
rect 1474 916 1477 933
rect 1482 923 1485 1016
rect 1490 1003 1493 1126
rect 1498 1106 1501 1126
rect 1498 1103 1509 1106
rect 1506 1046 1509 1103
rect 1498 1043 1509 1046
rect 1498 1023 1501 1043
rect 1490 916 1493 966
rect 1498 953 1501 1016
rect 1506 993 1509 1006
rect 1498 923 1501 946
rect 1506 933 1509 976
rect 1514 963 1517 1006
rect 1522 956 1525 1016
rect 1546 1013 1549 1126
rect 1554 1113 1557 1126
rect 1562 993 1565 1293
rect 1570 1203 1573 1216
rect 1586 1173 1589 1356
rect 1626 1246 1629 1373
rect 1642 1313 1645 1326
rect 1626 1243 1637 1246
rect 1578 1133 1581 1146
rect 1594 1133 1597 1206
rect 1602 1186 1605 1236
rect 1634 1223 1637 1243
rect 1642 1216 1645 1236
rect 1650 1233 1653 1406
rect 1662 1366 1665 1423
rect 1662 1363 1669 1366
rect 1666 1343 1669 1363
rect 1674 1336 1677 1416
rect 1698 1393 1701 1486
rect 1778 1483 1781 1756
rect 1714 1353 1717 1456
rect 1786 1446 1789 1846
rect 1810 1823 1813 1926
rect 1810 1793 1813 1816
rect 1794 1716 1797 1736
rect 1794 1713 1805 1716
rect 1802 1646 1805 1713
rect 1818 1653 1821 1933
rect 1826 1916 1829 2033
rect 1834 1973 1837 2113
rect 1834 1933 1837 1946
rect 1842 1933 1845 2106
rect 1866 2003 1869 2056
rect 1890 1993 1893 2166
rect 1906 2163 1909 2283
rect 1930 2216 1933 2326
rect 1970 2316 1973 2366
rect 1978 2323 1981 2346
rect 1970 2313 1981 2316
rect 1938 2223 1941 2236
rect 1914 2193 1917 2206
rect 1906 2123 1909 2146
rect 1858 1923 1861 1936
rect 1826 1913 1833 1916
rect 1830 1816 1833 1913
rect 1826 1813 1833 1816
rect 1826 1793 1829 1813
rect 1858 1736 1861 1836
rect 1866 1743 1869 1976
rect 1882 1926 1885 1946
rect 1906 1933 1909 1986
rect 1914 1943 1917 2026
rect 1874 1796 1877 1926
rect 1882 1923 1893 1926
rect 1890 1856 1893 1923
rect 1914 1876 1917 1936
rect 1922 1923 1925 2216
rect 1930 2213 1941 2216
rect 1938 2203 1941 2213
rect 1930 2116 1933 2196
rect 1954 2163 1957 2206
rect 1938 2133 1949 2136
rect 1930 2113 1937 2116
rect 1934 2046 1937 2113
rect 1946 2103 1949 2126
rect 1930 2043 1937 2046
rect 1930 2023 1933 2043
rect 1930 1933 1933 2016
rect 1946 1933 1949 1956
rect 1882 1853 1893 1856
rect 1906 1873 1917 1876
rect 1882 1833 1885 1853
rect 1882 1813 1885 1826
rect 1906 1813 1909 1873
rect 1922 1816 1925 1916
rect 1938 1913 1941 1926
rect 1954 1916 1957 2126
rect 1950 1913 1957 1916
rect 1950 1836 1953 1913
rect 1950 1833 1957 1836
rect 1914 1813 1933 1816
rect 1946 1806 1949 1816
rect 1954 1813 1957 1833
rect 1890 1803 1901 1806
rect 1874 1793 1881 1796
rect 1834 1696 1837 1736
rect 1858 1733 1869 1736
rect 1878 1726 1881 1793
rect 1842 1723 1861 1726
rect 1866 1716 1869 1726
rect 1878 1723 1885 1726
rect 1842 1713 1869 1716
rect 1834 1693 1845 1696
rect 1794 1643 1805 1646
rect 1794 1613 1797 1643
rect 1842 1636 1845 1693
rect 1874 1683 1877 1716
rect 1882 1693 1885 1723
rect 1834 1633 1845 1636
rect 1834 1613 1837 1633
rect 1890 1613 1893 1796
rect 1906 1773 1909 1806
rect 1906 1733 1909 1746
rect 1810 1593 1813 1606
rect 1802 1523 1805 1546
rect 1850 1533 1853 1596
rect 1898 1536 1901 1706
rect 1882 1533 1901 1536
rect 1906 1533 1909 1726
rect 1930 1696 1933 1766
rect 1938 1723 1941 1806
rect 1946 1803 1957 1806
rect 1954 1793 1957 1803
rect 1962 1786 1965 2156
rect 1970 2133 1973 2146
rect 1978 2103 1981 2313
rect 1994 2303 1997 2376
rect 2002 2363 2005 2406
rect 2026 2216 2029 2406
rect 2042 2403 2045 2413
rect 2058 2403 2061 2416
rect 2082 2413 2085 2473
rect 2074 2393 2077 2406
rect 2090 2386 2093 2483
rect 2098 2453 2101 2516
rect 2114 2473 2117 2536
rect 2146 2533 2165 2536
rect 2122 2453 2125 2526
rect 2138 2503 2141 2526
rect 2154 2503 2157 2526
rect 2162 2523 2165 2533
rect 2170 2506 2173 2566
rect 2166 2503 2173 2506
rect 2166 2436 2169 2503
rect 2162 2433 2169 2436
rect 2114 2393 2117 2416
rect 2162 2393 2165 2433
rect 2178 2403 2181 2506
rect 2186 2403 2189 2416
rect 2202 2403 2205 2526
rect 2210 2503 2213 2816
rect 2250 2813 2253 2883
rect 2314 2823 2317 2946
rect 2346 2933 2349 2946
rect 2234 2793 2237 2806
rect 2290 2793 2293 2816
rect 2338 2803 2341 2826
rect 2354 2803 2357 2816
rect 2218 2696 2221 2726
rect 2218 2693 2225 2696
rect 2222 2626 2225 2693
rect 2234 2643 2237 2736
rect 2282 2723 2285 2746
rect 2322 2733 2325 2746
rect 2274 2686 2277 2716
rect 2314 2713 2317 2726
rect 2330 2723 2341 2726
rect 2218 2623 2225 2626
rect 2258 2626 2261 2686
rect 2274 2683 2293 2686
rect 2258 2623 2269 2626
rect 2218 2603 2221 2623
rect 2242 2613 2261 2616
rect 2226 2573 2229 2606
rect 2242 2533 2245 2566
rect 2258 2563 2261 2606
rect 2226 2423 2229 2436
rect 2242 2413 2245 2526
rect 2250 2423 2253 2436
rect 2258 2426 2261 2536
rect 2266 2443 2269 2623
rect 2282 2613 2285 2636
rect 2274 2523 2277 2606
rect 2282 2583 2285 2606
rect 2290 2573 2293 2683
rect 2298 2566 2301 2656
rect 2306 2623 2309 2686
rect 2314 2616 2317 2706
rect 2322 2623 2325 2716
rect 2330 2703 2333 2723
rect 2306 2613 2317 2616
rect 2330 2613 2333 2646
rect 2306 2583 2309 2613
rect 2314 2573 2317 2606
rect 2338 2603 2341 2716
rect 2354 2713 2357 2736
rect 2362 2723 2365 2816
rect 2378 2803 2381 2926
rect 2426 2836 2429 2963
rect 2386 2823 2389 2836
rect 2418 2833 2429 2836
rect 2378 2723 2381 2746
rect 2410 2736 2413 2816
rect 2418 2803 2421 2833
rect 2434 2763 2437 2806
rect 2442 2803 2445 3040
rect 2642 2966 2645 3040
rect 2634 2963 2645 2966
rect 2522 2933 2525 2946
rect 2554 2933 2557 2946
rect 2450 2833 2461 2836
rect 2458 2823 2461 2833
rect 2466 2823 2493 2826
rect 2458 2793 2461 2816
rect 2466 2813 2469 2823
rect 2474 2803 2477 2816
rect 2498 2803 2501 2926
rect 2522 2813 2525 2826
rect 2578 2823 2581 2926
rect 2634 2856 2637 2963
rect 2666 2933 2669 2946
rect 2754 2933 2757 3040
rect 2626 2853 2637 2856
rect 2586 2823 2605 2826
rect 2610 2823 2613 2836
rect 2410 2733 2421 2736
rect 2346 2603 2349 2616
rect 2298 2563 2317 2566
rect 2274 2493 2277 2516
rect 2290 2466 2293 2556
rect 2314 2503 2317 2563
rect 2274 2463 2293 2466
rect 2258 2423 2269 2426
rect 2074 2383 2093 2386
rect 2058 2326 2061 2346
rect 2042 2303 2045 2326
rect 2058 2323 2065 2326
rect 2050 2243 2053 2286
rect 1986 2196 1989 2216
rect 1986 2193 1993 2196
rect 1990 2106 1993 2193
rect 1990 2103 1997 2106
rect 1970 1866 1973 2036
rect 1978 1883 1981 2026
rect 1986 1933 1989 2016
rect 1994 2003 1997 2103
rect 2002 2093 2005 2216
rect 2018 2213 2037 2216
rect 2042 2213 2045 2226
rect 2050 2213 2053 2236
rect 2062 2226 2065 2323
rect 2074 2283 2077 2383
rect 2090 2333 2093 2376
rect 2130 2336 2133 2366
rect 2122 2333 2133 2336
rect 2058 2223 2065 2226
rect 2018 2133 2021 2213
rect 2058 2203 2061 2223
rect 2066 2193 2069 2206
rect 2034 2133 2037 2156
rect 2074 2136 2077 2216
rect 2090 2203 2093 2306
rect 2098 2203 2101 2286
rect 2122 2276 2125 2333
rect 2138 2286 2141 2326
rect 2138 2283 2149 2286
rect 2122 2273 2133 2276
rect 2106 2223 2117 2226
rect 2122 2223 2125 2256
rect 2106 2213 2109 2223
rect 2010 2096 2013 2126
rect 2010 2093 2021 2096
rect 2018 2046 2021 2093
rect 2010 2043 2021 2046
rect 2010 2023 2013 2043
rect 1994 1933 1997 1946
rect 1986 1913 1989 1926
rect 1994 1923 2005 1926
rect 2002 1896 2005 1916
rect 1994 1893 2005 1896
rect 1970 1863 1977 1866
rect 1954 1783 1965 1786
rect 1954 1703 1957 1783
rect 1914 1603 1917 1626
rect 1922 1526 1925 1696
rect 1930 1693 1957 1696
rect 1938 1563 1941 1656
rect 1946 1593 1949 1606
rect 1938 1536 1941 1556
rect 1930 1533 1941 1536
rect 1786 1443 1797 1446
rect 1730 1413 1741 1416
rect 1754 1413 1765 1416
rect 1730 1403 1733 1413
rect 1754 1403 1757 1413
rect 1778 1393 1781 1406
rect 1794 1383 1797 1443
rect 1834 1426 1837 1486
rect 1866 1453 1869 1526
rect 1890 1523 1941 1526
rect 1826 1423 1837 1426
rect 1626 1213 1645 1216
rect 1610 1193 1621 1196
rect 1626 1193 1629 1206
rect 1602 1183 1613 1186
rect 1586 1023 1589 1126
rect 1586 1003 1589 1016
rect 1514 953 1525 956
rect 1474 913 1485 916
rect 1490 913 1501 916
rect 1402 843 1413 846
rect 1410 813 1413 843
rect 1418 813 1421 846
rect 1442 843 1453 846
rect 1378 756 1381 806
rect 1386 803 1405 806
rect 1426 756 1429 826
rect 1434 766 1437 826
rect 1450 803 1453 843
rect 1458 823 1469 826
rect 1458 803 1461 816
rect 1466 813 1469 823
rect 1474 813 1477 896
rect 1482 813 1485 913
rect 1498 836 1501 913
rect 1514 846 1517 953
rect 1522 913 1525 936
rect 1554 933 1557 946
rect 1578 933 1581 956
rect 1530 913 1557 916
rect 1514 843 1525 846
rect 1498 833 1509 836
rect 1506 813 1509 833
rect 1522 806 1525 843
rect 1474 803 1485 806
rect 1498 793 1501 806
rect 1514 803 1525 806
rect 1434 763 1469 766
rect 1370 753 1381 756
rect 1298 716 1301 736
rect 1306 723 1309 746
rect 1318 743 1325 746
rect 1322 726 1325 743
rect 1322 723 1329 726
rect 1370 723 1373 753
rect 1394 733 1397 756
rect 1418 753 1429 756
rect 1274 713 1285 716
rect 1298 713 1317 716
rect 1194 573 1213 576
rect 1186 503 1189 526
rect 1194 496 1197 536
rect 1186 493 1197 496
rect 1106 373 1109 406
rect 1130 393 1133 416
rect 994 163 997 206
rect 1010 166 1013 206
rect 1034 193 1037 216
rect 1090 213 1093 356
rect 1114 323 1117 346
rect 1106 213 1109 226
rect 1114 213 1125 216
rect 1130 213 1133 236
rect 1146 213 1149 226
rect 1122 193 1125 213
rect 1002 163 1013 166
rect 1002 133 1005 163
rect 1026 123 1029 146
rect 1106 133 1109 186
rect 1082 113 1085 126
rect 1138 123 1141 206
rect 1154 143 1157 206
rect 1162 183 1165 376
rect 1178 323 1181 406
rect 1186 333 1189 493
rect 1202 483 1205 526
rect 1210 406 1213 573
rect 1218 533 1221 596
rect 1234 593 1245 596
rect 1250 663 1261 666
rect 1250 593 1253 663
rect 1282 603 1285 713
rect 1290 613 1293 626
rect 1314 613 1317 713
rect 1326 626 1329 723
rect 1322 623 1329 626
rect 1338 623 1341 636
rect 1234 493 1237 593
rect 1290 566 1293 596
rect 1290 563 1301 566
rect 1282 523 1285 546
rect 1298 513 1301 563
rect 1306 533 1309 606
rect 1322 603 1325 623
rect 1314 523 1317 596
rect 1338 593 1341 606
rect 1346 573 1349 616
rect 1354 613 1357 626
rect 1362 613 1365 656
rect 1370 603 1373 626
rect 1386 613 1389 686
rect 1418 683 1421 753
rect 1434 703 1437 736
rect 1466 666 1469 763
rect 1522 743 1525 766
rect 1530 736 1533 913
rect 1562 903 1565 926
rect 1594 923 1597 1066
rect 1602 1013 1605 1156
rect 1610 933 1613 1183
rect 1618 1153 1621 1193
rect 1642 1176 1645 1196
rect 1634 1173 1645 1176
rect 1618 1103 1621 1126
rect 1634 1066 1637 1173
rect 1650 1133 1653 1216
rect 1658 1143 1661 1226
rect 1666 1216 1669 1336
rect 1674 1333 1693 1336
rect 1714 1333 1717 1346
rect 1730 1333 1733 1366
rect 1754 1336 1757 1356
rect 1754 1333 1765 1336
rect 1674 1223 1677 1236
rect 1666 1213 1677 1216
rect 1634 1063 1645 1066
rect 1634 933 1637 1046
rect 1642 993 1645 1063
rect 1650 1053 1653 1126
rect 1674 1123 1677 1213
rect 1682 1186 1685 1326
rect 1690 1226 1693 1316
rect 1714 1303 1717 1326
rect 1762 1256 1765 1333
rect 1778 1313 1781 1326
rect 1746 1253 1765 1256
rect 1746 1236 1749 1253
rect 1698 1233 1717 1236
rect 1714 1226 1717 1233
rect 1742 1233 1749 1236
rect 1690 1223 1709 1226
rect 1714 1223 1733 1226
rect 1690 1193 1693 1216
rect 1714 1203 1717 1223
rect 1682 1183 1709 1186
rect 1674 1023 1677 1036
rect 1658 996 1661 1016
rect 1682 1013 1685 1136
rect 1690 1023 1693 1146
rect 1706 1106 1709 1183
rect 1702 1103 1709 1106
rect 1702 1036 1705 1103
rect 1722 1086 1725 1216
rect 1730 1213 1733 1223
rect 1742 1176 1745 1233
rect 1742 1173 1749 1176
rect 1746 1126 1749 1173
rect 1762 1133 1765 1216
rect 1810 1183 1813 1396
rect 1826 1356 1829 1423
rect 1842 1376 1845 1416
rect 1842 1373 1853 1376
rect 1826 1353 1837 1356
rect 1826 1213 1829 1326
rect 1826 1193 1829 1206
rect 1802 1146 1805 1166
rect 1834 1163 1837 1353
rect 1850 1333 1853 1373
rect 1866 1333 1869 1406
rect 1890 1403 1893 1416
rect 1882 1333 1885 1346
rect 1842 1323 1853 1326
rect 1842 1203 1845 1316
rect 1858 1303 1861 1326
rect 1802 1143 1813 1146
rect 1746 1123 1757 1126
rect 1698 1033 1705 1036
rect 1714 1083 1725 1086
rect 1650 993 1661 996
rect 1578 846 1581 916
rect 1570 843 1581 846
rect 1522 733 1533 736
rect 1538 726 1541 836
rect 1554 793 1557 816
rect 1570 776 1573 843
rect 1610 833 1613 916
rect 1618 893 1621 926
rect 1650 923 1653 993
rect 1666 966 1669 1006
rect 1682 976 1685 1006
rect 1690 993 1693 1016
rect 1698 1003 1701 1033
rect 1714 1023 1717 1083
rect 1722 1023 1725 1056
rect 1706 996 1709 1016
rect 1698 993 1709 996
rect 1682 973 1689 976
rect 1666 963 1677 966
rect 1674 933 1677 963
rect 1666 883 1669 916
rect 1674 863 1677 926
rect 1686 906 1689 973
rect 1698 923 1701 993
rect 1714 923 1717 936
rect 1722 923 1725 996
rect 1730 933 1733 1036
rect 1738 1023 1741 1036
rect 1746 1023 1749 1116
rect 1754 1106 1757 1123
rect 1754 1103 1761 1106
rect 1758 1016 1761 1103
rect 1754 1013 1761 1016
rect 1754 926 1757 1013
rect 1778 993 1781 1136
rect 1810 1096 1813 1143
rect 1826 1123 1829 1136
rect 1802 1093 1813 1096
rect 1802 996 1805 1093
rect 1850 1026 1853 1236
rect 1858 1196 1861 1206
rect 1866 1203 1869 1216
rect 1874 1196 1877 1216
rect 1858 1193 1877 1196
rect 1874 1066 1877 1193
rect 1882 1133 1885 1206
rect 1874 1063 1881 1066
rect 1846 1023 1853 1026
rect 1794 993 1805 996
rect 1746 923 1757 926
rect 1682 903 1689 906
rect 1682 883 1685 903
rect 1434 663 1469 666
rect 1394 613 1397 626
rect 1386 563 1389 596
rect 1322 533 1325 556
rect 1330 526 1333 536
rect 1346 533 1357 536
rect 1330 523 1349 526
rect 1354 523 1357 533
rect 1370 526 1373 536
rect 1394 533 1397 606
rect 1410 543 1413 606
rect 1370 523 1381 526
rect 1218 413 1253 416
rect 1194 373 1197 406
rect 1210 403 1229 406
rect 1202 286 1205 336
rect 1210 323 1213 336
rect 1218 333 1221 346
rect 1202 283 1213 286
rect 1170 193 1173 206
rect 1178 203 1181 216
rect 1194 213 1197 226
rect 1186 133 1189 206
rect 1202 173 1205 206
rect 1210 193 1213 283
rect 1218 213 1221 276
rect 1226 226 1229 403
rect 1234 333 1237 406
rect 1258 366 1261 496
rect 1266 403 1269 416
rect 1282 373 1285 486
rect 1330 413 1333 516
rect 1346 513 1373 516
rect 1378 413 1381 523
rect 1394 513 1397 526
rect 1418 523 1421 616
rect 1434 613 1437 663
rect 1458 613 1461 656
rect 1482 626 1485 726
rect 1514 646 1517 726
rect 1506 643 1517 646
rect 1530 723 1541 726
rect 1466 616 1469 626
rect 1482 623 1501 626
rect 1466 613 1477 616
rect 1426 543 1429 606
rect 1434 583 1437 596
rect 1458 593 1461 606
rect 1466 563 1469 606
rect 1426 523 1429 536
rect 1474 533 1477 613
rect 1482 593 1485 616
rect 1490 553 1493 606
rect 1498 563 1501 623
rect 1506 603 1509 643
rect 1530 636 1533 723
rect 1546 706 1549 726
rect 1554 723 1557 776
rect 1570 773 1581 776
rect 1578 756 1581 773
rect 1578 753 1589 756
rect 1602 753 1605 806
rect 1626 793 1629 806
rect 1658 793 1661 816
rect 1698 766 1701 916
rect 1714 883 1717 916
rect 1746 913 1749 923
rect 1754 883 1757 916
rect 1762 913 1765 946
rect 1770 933 1781 936
rect 1778 913 1781 926
rect 1690 763 1701 766
rect 1570 743 1581 746
rect 1562 733 1573 736
rect 1586 726 1589 753
rect 1570 723 1589 726
rect 1514 633 1533 636
rect 1538 703 1549 706
rect 1514 613 1517 633
rect 1514 593 1517 606
rect 1530 603 1533 626
rect 1538 613 1541 703
rect 1554 616 1557 716
rect 1554 613 1565 616
rect 1570 613 1573 723
rect 1594 713 1597 726
rect 1610 636 1613 736
rect 1634 713 1637 726
rect 1690 716 1693 763
rect 1706 723 1709 736
rect 1714 733 1717 816
rect 1722 813 1725 866
rect 1690 713 1701 716
rect 1730 713 1733 816
rect 1738 793 1741 806
rect 1746 783 1749 846
rect 1754 823 1765 826
rect 1610 633 1621 636
rect 1578 613 1581 626
rect 1602 616 1605 626
rect 1594 613 1605 616
rect 1434 513 1445 516
rect 1394 486 1397 506
rect 1394 483 1405 486
rect 1402 426 1405 483
rect 1442 433 1445 513
rect 1394 423 1405 426
rect 1298 393 1301 406
rect 1250 363 1261 366
rect 1250 333 1253 363
rect 1386 356 1389 406
rect 1394 403 1397 423
rect 1426 406 1429 426
rect 1418 403 1429 406
rect 1378 346 1381 356
rect 1386 353 1397 356
rect 1234 313 1237 326
rect 1250 286 1253 326
rect 1274 323 1277 346
rect 1370 343 1389 346
rect 1338 333 1357 336
rect 1338 323 1349 326
rect 1338 293 1341 323
rect 1250 283 1261 286
rect 1226 223 1237 226
rect 1234 213 1237 223
rect 1242 213 1245 226
rect 1226 193 1229 206
rect 1210 133 1213 166
rect 1218 123 1221 146
rect 1242 133 1245 156
rect 1258 153 1261 283
rect 1282 193 1285 216
rect 1346 213 1349 316
rect 1354 303 1357 333
rect 1370 326 1373 343
rect 1366 323 1373 326
rect 1378 323 1381 336
rect 1394 326 1397 353
rect 1434 346 1437 406
rect 1386 323 1397 326
rect 1366 236 1369 323
rect 1366 233 1373 236
rect 1354 213 1357 226
rect 1370 213 1373 233
rect 1266 123 1269 136
rect 1330 123 1333 156
rect 1338 123 1341 176
rect 1346 113 1349 206
rect 1362 163 1365 206
rect 1370 146 1373 186
rect 1362 143 1373 146
rect 1378 143 1381 296
rect 1386 206 1389 323
rect 1394 303 1397 316
rect 1402 313 1405 326
rect 1410 303 1413 346
rect 1434 343 1445 346
rect 1418 233 1421 326
rect 1426 253 1429 336
rect 1394 213 1397 226
rect 1386 203 1397 206
rect 1378 123 1381 136
rect 1386 113 1389 126
rect 1394 106 1397 146
rect 1402 123 1405 226
rect 1426 213 1429 226
rect 1410 166 1413 206
rect 1410 163 1421 166
rect 1418 133 1421 163
rect 1434 126 1437 326
rect 1442 293 1445 343
rect 1450 333 1453 526
rect 1458 423 1461 526
rect 1466 523 1477 526
rect 1474 476 1477 516
rect 1466 473 1477 476
rect 1466 406 1469 473
rect 1474 423 1477 436
rect 1482 423 1485 546
rect 1490 526 1493 536
rect 1490 523 1525 526
rect 1490 513 1493 523
rect 1474 413 1501 416
rect 1458 343 1461 406
rect 1466 403 1477 406
rect 1450 313 1453 326
rect 1458 266 1461 316
rect 1466 313 1469 326
rect 1450 263 1461 266
rect 1442 213 1445 226
rect 1442 133 1445 156
rect 1450 133 1453 263
rect 1458 223 1461 256
rect 1466 216 1469 306
rect 1474 243 1477 403
rect 1506 356 1509 426
rect 1498 353 1509 356
rect 1482 333 1493 336
rect 1482 313 1485 333
rect 1498 326 1501 353
rect 1514 346 1517 406
rect 1490 323 1501 326
rect 1506 343 1517 346
rect 1506 323 1509 343
rect 1522 336 1525 436
rect 1530 413 1533 446
rect 1546 426 1549 536
rect 1554 513 1557 606
rect 1562 586 1565 613
rect 1570 593 1573 606
rect 1578 586 1581 606
rect 1562 583 1573 586
rect 1578 583 1589 586
rect 1562 533 1565 546
rect 1562 503 1565 526
rect 1570 496 1573 583
rect 1578 533 1581 556
rect 1586 533 1589 583
rect 1578 513 1581 526
rect 1594 516 1597 613
rect 1602 593 1605 606
rect 1590 513 1597 516
rect 1562 493 1573 496
rect 1538 413 1541 426
rect 1546 423 1557 426
rect 1514 333 1525 336
rect 1538 323 1541 406
rect 1546 323 1549 416
rect 1466 213 1477 216
rect 1466 186 1469 206
rect 1458 183 1469 186
rect 1458 133 1461 183
rect 1434 123 1445 126
rect 1402 113 1413 116
rect 1442 113 1453 116
rect 1458 113 1461 126
rect 1466 123 1469 136
rect 1474 113 1477 213
rect 1482 183 1485 226
rect 1490 193 1493 323
rect 1498 203 1501 246
rect 1506 213 1509 226
rect 1514 216 1517 276
rect 1530 233 1533 316
rect 1538 243 1541 316
rect 1554 313 1557 423
rect 1562 403 1565 493
rect 1590 446 1593 513
rect 1590 443 1597 446
rect 1522 223 1533 226
rect 1514 213 1525 216
rect 1538 136 1541 236
rect 1546 226 1549 236
rect 1546 223 1557 226
rect 1546 173 1549 216
rect 1482 113 1485 136
rect 1514 133 1541 136
rect 1554 113 1557 223
rect 1562 203 1565 346
rect 1570 336 1573 436
rect 1586 413 1589 426
rect 1594 413 1597 443
rect 1594 356 1597 406
rect 1602 403 1605 556
rect 1618 553 1621 633
rect 1642 593 1645 616
rect 1610 403 1613 506
rect 1618 403 1621 516
rect 1634 513 1637 536
rect 1650 533 1653 556
rect 1674 513 1677 526
rect 1690 506 1693 526
rect 1686 503 1693 506
rect 1626 423 1629 446
rect 1686 436 1689 503
rect 1634 423 1637 436
rect 1686 433 1693 436
rect 1626 403 1629 416
rect 1634 406 1637 416
rect 1634 403 1661 406
rect 1586 353 1597 356
rect 1570 333 1581 336
rect 1570 303 1573 326
rect 1578 273 1581 333
rect 1586 233 1589 353
rect 1594 343 1613 346
rect 1610 333 1613 343
rect 1618 333 1637 336
rect 1594 316 1597 326
rect 1602 323 1613 326
rect 1618 323 1621 333
rect 1594 313 1621 316
rect 1626 313 1629 326
rect 1634 313 1637 333
rect 1594 233 1597 306
rect 1578 223 1589 226
rect 1578 216 1581 223
rect 1570 213 1581 216
rect 1562 123 1565 196
rect 1586 133 1589 216
rect 1594 173 1597 216
rect 1602 196 1605 236
rect 1610 213 1613 226
rect 1642 223 1645 336
rect 1650 273 1653 326
rect 1666 313 1669 406
rect 1674 396 1677 416
rect 1690 413 1693 433
rect 1674 393 1685 396
rect 1682 336 1685 393
rect 1674 333 1685 336
rect 1674 313 1677 333
rect 1658 256 1661 306
rect 1658 253 1669 256
rect 1634 213 1653 216
rect 1666 213 1669 253
rect 1634 203 1637 213
rect 1602 193 1613 196
rect 1642 193 1645 206
rect 866 103 877 106
rect 1394 103 1413 106
rect 1586 103 1589 116
rect 1594 113 1597 126
rect 1602 123 1605 186
rect 1610 103 1613 193
rect 1618 103 1621 116
rect -622 -659 -56 -654
rect -43 3 0 8
rect -865 -733 -859 -727
rect -862 -739 -859 -733
rect -852 -748 -846 -737
rect -622 -743 -617 -659
rect -43 -676 -38 3
rect 1698 0 1701 713
rect 1706 606 1709 616
rect 1714 613 1717 626
rect 1706 603 1725 606
rect 1738 603 1741 776
rect 1754 753 1757 806
rect 1762 766 1765 823
rect 1770 773 1773 906
rect 1786 866 1789 936
rect 1794 903 1797 993
rect 1810 933 1813 1016
rect 1802 913 1805 926
rect 1778 863 1789 866
rect 1778 813 1781 863
rect 1794 823 1813 826
rect 1794 813 1797 823
rect 1802 806 1805 816
rect 1786 803 1805 806
rect 1810 793 1813 823
rect 1818 773 1821 946
rect 1846 936 1849 1023
rect 1846 933 1853 936
rect 1858 933 1861 1016
rect 1866 1013 1869 1056
rect 1842 896 1845 916
rect 1838 893 1845 896
rect 1838 776 1841 893
rect 1838 773 1845 776
rect 1762 763 1773 766
rect 1770 746 1773 763
rect 1754 733 1757 746
rect 1770 743 1789 746
rect 1754 583 1757 726
rect 1786 696 1789 743
rect 1802 723 1805 746
rect 1842 733 1845 773
rect 1834 723 1845 726
rect 1850 723 1853 933
rect 1866 923 1869 1006
rect 1878 996 1881 1063
rect 1878 993 1885 996
rect 1874 913 1877 926
rect 1882 923 1885 993
rect 1890 913 1893 1216
rect 1898 1213 1901 1226
rect 1906 1213 1909 1516
rect 1938 1513 1941 1523
rect 1946 1496 1949 1546
rect 1938 1493 1949 1496
rect 1938 1363 1941 1493
rect 1954 1443 1957 1693
rect 1974 1686 1977 1863
rect 1994 1836 1997 1893
rect 1994 1833 2005 1836
rect 2002 1813 2005 1833
rect 2010 1813 2013 1986
rect 2026 1926 2029 2016
rect 2034 1983 2037 2006
rect 2018 1923 2029 1926
rect 1986 1723 1989 1806
rect 1994 1753 1997 1806
rect 2010 1766 2013 1806
rect 2018 1773 2021 1906
rect 2042 1876 2045 2016
rect 2058 2003 2061 2136
rect 2070 2133 2077 2136
rect 2070 2006 2073 2133
rect 2082 2016 2085 2126
rect 2114 2116 2117 2216
rect 2130 2136 2133 2273
rect 2138 2203 2141 2276
rect 2146 2203 2149 2283
rect 2170 2273 2173 2386
rect 2194 2333 2197 2376
rect 2210 2343 2213 2406
rect 2226 2383 2229 2406
rect 2250 2403 2253 2416
rect 2266 2396 2269 2423
rect 2274 2403 2277 2463
rect 2314 2413 2317 2436
rect 2266 2393 2277 2396
rect 2178 2223 2181 2236
rect 2162 2186 2165 2216
rect 2154 2183 2165 2186
rect 2122 2133 2141 2136
rect 2122 2123 2125 2133
rect 2114 2113 2125 2116
rect 2090 2023 2093 2086
rect 2130 2083 2133 2126
rect 2154 2026 2157 2183
rect 2146 2023 2157 2026
rect 2082 2013 2093 2016
rect 2070 2003 2077 2006
rect 2090 2003 2093 2013
rect 2066 1923 2069 1946
rect 2074 1916 2077 2003
rect 2106 1976 2109 2006
rect 2106 1973 2117 1976
rect 2038 1873 2045 1876
rect 2066 1913 2077 1916
rect 2026 1813 2029 1826
rect 2038 1816 2041 1873
rect 2034 1813 2041 1816
rect 2050 1813 2053 1866
rect 2026 1793 2029 1806
rect 2010 1763 2029 1766
rect 2002 1733 2005 1746
rect 2026 1723 2029 1763
rect 2034 1716 2037 1813
rect 2042 1803 2053 1806
rect 1970 1683 1977 1686
rect 1962 1613 1965 1626
rect 1962 1513 1965 1526
rect 1970 1503 1973 1683
rect 1986 1603 1989 1716
rect 2026 1713 2037 1716
rect 2042 1716 2045 1776
rect 2050 1723 2053 1803
rect 2058 1783 2061 1836
rect 2066 1813 2069 1913
rect 2090 1873 2093 1946
rect 2042 1713 2053 1716
rect 1994 1613 1997 1626
rect 1994 1603 2013 1606
rect 2018 1603 2021 1636
rect 2026 1613 2029 1713
rect 1978 1523 1981 1536
rect 1994 1533 1997 1603
rect 2018 1546 2021 1566
rect 2018 1543 2025 1546
rect 2022 1476 2025 1543
rect 2034 1523 2037 1606
rect 2042 1603 2045 1616
rect 2018 1473 2025 1476
rect 2018 1456 2021 1473
rect 2010 1453 2021 1456
rect 2042 1456 2045 1576
rect 2050 1566 2053 1713
rect 2066 1706 2069 1806
rect 2074 1756 2077 1806
rect 2074 1753 2085 1756
rect 2082 1723 2085 1753
rect 2090 1743 2093 1816
rect 2114 1813 2117 1973
rect 2130 1933 2133 2016
rect 2146 1996 2149 2023
rect 2154 2003 2157 2016
rect 2146 1993 2157 1996
rect 2090 1723 2093 1736
rect 2098 1706 2101 1766
rect 2122 1763 2125 1826
rect 2130 1806 2133 1926
rect 2138 1863 2141 1926
rect 2146 1856 2149 1936
rect 2154 1926 2157 1993
rect 2170 1946 2173 2206
rect 2194 2193 2197 2206
rect 2178 2106 2181 2126
rect 2202 2113 2205 2216
rect 2210 2183 2213 2206
rect 2210 2133 2213 2146
rect 2218 2106 2221 2216
rect 2234 2203 2237 2326
rect 2242 2213 2245 2226
rect 2274 2213 2277 2393
rect 2282 2363 2285 2406
rect 2322 2403 2325 2526
rect 2354 2523 2357 2636
rect 2362 2613 2365 2626
rect 2370 2613 2373 2696
rect 2402 2656 2405 2726
rect 2394 2653 2405 2656
rect 2386 2623 2389 2636
rect 2394 2616 2397 2653
rect 2418 2646 2421 2733
rect 2458 2666 2461 2766
rect 2522 2756 2525 2806
rect 2522 2753 2533 2756
rect 2466 2723 2469 2736
rect 2450 2663 2461 2666
rect 2410 2643 2421 2646
rect 2386 2613 2397 2616
rect 2362 2413 2365 2566
rect 2370 2523 2373 2606
rect 2378 2533 2381 2606
rect 2386 2603 2389 2613
rect 2402 2583 2405 2616
rect 2410 2603 2413 2643
rect 2418 2593 2421 2626
rect 2426 2566 2429 2616
rect 2434 2613 2437 2646
rect 2442 2596 2445 2606
rect 2450 2603 2453 2663
rect 2458 2596 2461 2616
rect 2442 2593 2461 2596
rect 2426 2563 2453 2566
rect 2418 2533 2421 2556
rect 2370 2403 2373 2506
rect 2386 2483 2389 2526
rect 2402 2436 2405 2526
rect 2442 2486 2445 2526
rect 2438 2483 2445 2486
rect 2394 2433 2405 2436
rect 2386 2386 2389 2406
rect 2382 2383 2389 2386
rect 2290 2333 2293 2376
rect 2258 2203 2269 2206
rect 2282 2186 2285 2216
rect 2274 2183 2285 2186
rect 2178 2103 2189 2106
rect 2186 2026 2189 2103
rect 2178 2023 2189 2026
rect 2202 2103 2221 2106
rect 2178 1973 2181 2023
rect 2162 1933 2165 1946
rect 2170 1943 2181 1946
rect 2154 1923 2165 1926
rect 2162 1913 2165 1923
rect 2170 1903 2173 1936
rect 2178 1933 2181 1943
rect 2186 1933 2189 2006
rect 2202 1956 2205 2103
rect 2234 2056 2237 2156
rect 2258 2123 2261 2146
rect 2274 2076 2277 2183
rect 2290 2173 2293 2206
rect 2314 2203 2317 2326
rect 2314 2123 2317 2196
rect 2322 2143 2325 2226
rect 2338 2203 2341 2306
rect 2370 2303 2373 2326
rect 2382 2236 2385 2383
rect 2394 2246 2397 2433
rect 2418 2426 2421 2446
rect 2402 2336 2405 2426
rect 2414 2423 2421 2426
rect 2414 2356 2417 2423
rect 2414 2353 2421 2356
rect 2402 2333 2413 2336
rect 2410 2293 2413 2333
rect 2394 2243 2401 2246
rect 2382 2233 2389 2236
rect 2330 2136 2333 2176
rect 2354 2153 2357 2216
rect 2322 2133 2333 2136
rect 2274 2073 2285 2076
rect 2218 2053 2237 2056
rect 2282 2056 2285 2073
rect 2282 2053 2293 2056
rect 2218 2003 2221 2053
rect 2194 1953 2205 1956
rect 2138 1853 2149 1856
rect 2138 1813 2141 1853
rect 2154 1846 2157 1896
rect 2178 1863 2181 1926
rect 2194 1923 2197 1953
rect 2154 1843 2165 1846
rect 2130 1803 2141 1806
rect 2066 1703 2077 1706
rect 2074 1626 2077 1703
rect 2058 1613 2061 1626
rect 2066 1623 2077 1626
rect 2090 1703 2101 1706
rect 2090 1626 2093 1703
rect 2106 1633 2109 1716
rect 2090 1623 2101 1626
rect 2050 1563 2061 1566
rect 2042 1453 2049 1456
rect 1954 1423 1957 1436
rect 1954 1393 1957 1406
rect 1970 1386 1973 1406
rect 1994 1393 1997 1416
rect 1946 1383 1973 1386
rect 1946 1366 1949 1383
rect 2010 1376 2013 1453
rect 2010 1373 2021 1376
rect 1946 1363 1953 1366
rect 1898 1133 1901 1206
rect 1906 1183 1909 1206
rect 1914 1193 1917 1326
rect 1922 1216 1925 1326
rect 1930 1223 1933 1316
rect 1950 1286 1953 1363
rect 1962 1316 1965 1366
rect 2018 1353 2021 1373
rect 2034 1366 2037 1446
rect 2046 1366 2049 1453
rect 2030 1363 2037 1366
rect 2042 1363 2049 1366
rect 2058 1366 2061 1563
rect 2066 1506 2069 1623
rect 2074 1523 2077 1606
rect 2098 1573 2101 1623
rect 2122 1603 2125 1726
rect 2090 1533 2093 1566
rect 2130 1523 2133 1606
rect 2138 1543 2141 1803
rect 2162 1776 2165 1843
rect 2186 1813 2189 1916
rect 2154 1773 2165 1776
rect 2154 1756 2157 1773
rect 2150 1753 2157 1756
rect 2150 1706 2153 1753
rect 2170 1733 2173 1746
rect 2194 1733 2197 1876
rect 2202 1833 2205 1946
rect 2210 1823 2213 1936
rect 2218 1863 2221 1926
rect 2226 1856 2229 1936
rect 2242 1933 2245 1946
rect 2250 1916 2253 2046
rect 2258 1976 2261 2026
rect 2266 1993 2269 2016
rect 2290 1986 2293 2053
rect 2322 2013 2325 2126
rect 2330 2013 2341 2016
rect 2282 1983 2293 1986
rect 2258 1973 2265 1976
rect 2246 1913 2253 1916
rect 2226 1853 2237 1856
rect 2234 1813 2237 1853
rect 2150 1703 2157 1706
rect 2146 1603 2149 1636
rect 2066 1503 2085 1506
rect 2066 1393 2069 1416
rect 2074 1413 2077 1436
rect 2082 1413 2085 1503
rect 2154 1483 2157 1703
rect 2162 1583 2165 1616
rect 2058 1363 2077 1366
rect 1970 1333 1989 1336
rect 1970 1323 1973 1333
rect 1962 1313 1973 1316
rect 1978 1313 1981 1326
rect 1946 1283 1953 1286
rect 1922 1213 1933 1216
rect 1898 1096 1901 1116
rect 1898 1093 1909 1096
rect 1906 1046 1909 1093
rect 1898 1043 1909 1046
rect 1898 1003 1901 1043
rect 1922 1033 1925 1206
rect 1930 1113 1933 1196
rect 1906 1013 1909 1026
rect 1922 1003 1925 1026
rect 1922 933 1925 996
rect 1946 993 1949 1283
rect 1970 1223 1973 1313
rect 1970 1196 1973 1216
rect 1962 1193 1973 1196
rect 1962 1133 1965 1193
rect 1978 1176 1981 1306
rect 1986 1263 1989 1333
rect 2002 1293 2005 1346
rect 2030 1266 2033 1363
rect 2042 1313 2045 1363
rect 2050 1323 2053 1346
rect 2030 1263 2037 1266
rect 2034 1243 2037 1263
rect 1974 1173 1981 1176
rect 1858 733 1861 816
rect 1866 723 1869 796
rect 1874 746 1877 776
rect 1882 756 1885 816
rect 1898 813 1901 916
rect 1946 886 1949 926
rect 1942 883 1949 886
rect 1930 826 1933 846
rect 1922 823 1933 826
rect 1898 763 1901 806
rect 1882 753 1901 756
rect 1874 743 1893 746
rect 1874 733 1877 743
rect 1874 713 1877 726
rect 1882 703 1885 736
rect 1778 693 1789 696
rect 1762 593 1765 606
rect 1730 523 1733 546
rect 1738 523 1741 536
rect 1770 516 1773 616
rect 1778 613 1781 693
rect 1890 683 1893 743
rect 1898 676 1901 753
rect 1906 733 1909 746
rect 1922 736 1925 823
rect 1942 816 1945 883
rect 1930 813 1945 816
rect 1930 803 1933 813
rect 1914 723 1917 736
rect 1922 733 1933 736
rect 1882 673 1901 676
rect 1786 603 1789 626
rect 1802 603 1805 616
rect 1826 593 1829 616
rect 1778 523 1781 556
rect 1762 513 1773 516
rect 1762 466 1765 513
rect 1762 463 1773 466
rect 1746 413 1749 426
rect 1770 413 1773 463
rect 1786 423 1789 536
rect 1794 433 1797 576
rect 1802 493 1805 586
rect 1834 526 1837 536
rect 1842 533 1845 616
rect 1810 506 1813 526
rect 1834 523 1861 526
rect 1858 513 1861 523
rect 1882 506 1885 673
rect 1898 646 1901 666
rect 1894 643 1901 646
rect 1894 546 1897 643
rect 1906 546 1909 626
rect 1914 603 1917 716
rect 1930 713 1933 733
rect 1938 713 1941 766
rect 1938 656 1941 706
rect 1946 663 1949 736
rect 1954 706 1957 1026
rect 1962 976 1965 1116
rect 1974 1076 1977 1173
rect 1974 1073 1981 1076
rect 1978 1056 1981 1073
rect 1986 1066 1989 1226
rect 1994 1133 1997 1146
rect 1986 1063 1997 1066
rect 1978 1053 1989 1056
rect 1970 993 1973 1016
rect 1986 1013 1989 1053
rect 1994 996 1997 1063
rect 1990 993 1997 996
rect 1962 973 1969 976
rect 1966 866 1969 973
rect 1990 886 1993 993
rect 2002 933 2005 1036
rect 1962 863 1969 866
rect 1978 883 1993 886
rect 1962 843 1965 863
rect 1970 803 1973 836
rect 1978 823 1981 883
rect 2002 833 2005 926
rect 1986 793 1989 816
rect 1994 803 1997 826
rect 2010 803 2013 1166
rect 2026 1143 2029 1216
rect 2042 1163 2045 1296
rect 2066 1203 2069 1356
rect 2058 1123 2061 1146
rect 2018 963 2021 1066
rect 2026 933 2029 1026
rect 2034 966 2037 1016
rect 2042 1013 2045 1026
rect 2058 1013 2069 1016
rect 2050 993 2053 1006
rect 2058 1003 2069 1006
rect 2034 963 2053 966
rect 2050 923 2053 963
rect 1978 723 1981 736
rect 1986 733 1989 786
rect 2010 713 2013 796
rect 1954 703 1965 706
rect 1938 653 1949 656
rect 1938 623 1941 636
rect 1946 623 1949 653
rect 1962 646 1965 703
rect 1954 643 1965 646
rect 1922 553 1925 616
rect 1938 556 1941 616
rect 1946 593 1949 606
rect 1930 553 1941 556
rect 1894 543 1901 546
rect 1906 543 1925 546
rect 1890 513 1893 526
rect 1810 503 1821 506
rect 1882 503 1893 506
rect 1818 436 1821 503
rect 1810 433 1821 436
rect 1714 333 1717 376
rect 1738 323 1741 396
rect 1770 383 1773 406
rect 1786 393 1789 406
rect 1810 373 1813 433
rect 1818 403 1821 416
rect 1842 393 1845 406
rect 1850 403 1853 416
rect 1866 413 1869 456
rect 1786 316 1789 356
rect 1794 323 1797 336
rect 1818 333 1821 366
rect 1850 333 1853 346
rect 1858 333 1861 406
rect 1874 343 1877 496
rect 1786 313 1797 316
rect 1794 166 1797 313
rect 1858 303 1861 326
rect 1866 256 1869 336
rect 1882 333 1885 396
rect 1890 363 1893 503
rect 1898 493 1901 543
rect 1906 353 1909 536
rect 1914 476 1917 536
rect 1922 523 1925 543
rect 1930 526 1933 553
rect 1938 533 1941 546
rect 1954 533 1957 643
rect 1962 563 1965 606
rect 1978 566 1981 616
rect 2002 593 2005 616
rect 1978 563 1997 566
rect 1930 523 1941 526
rect 1978 523 1981 546
rect 1938 513 1941 523
rect 1994 516 1997 563
rect 1986 513 1997 516
rect 1914 473 1925 476
rect 1922 396 1925 473
rect 1914 393 1925 396
rect 1914 373 1917 393
rect 1946 363 1949 406
rect 1970 396 1973 446
rect 1962 393 1973 396
rect 1890 333 1909 336
rect 1842 253 1869 256
rect 1786 163 1797 166
rect 1786 133 1789 163
rect 1834 123 1837 216
rect 1842 213 1845 253
rect 1882 213 1885 226
rect 1890 213 1893 333
rect 1898 316 1901 326
rect 1906 323 1909 333
rect 1898 313 1909 316
rect 1898 213 1901 226
rect 1906 213 1909 313
rect 1914 213 1917 336
rect 1922 306 1925 336
rect 1930 333 1933 346
rect 1954 326 1957 346
rect 1946 323 1957 326
rect 1922 303 1933 306
rect 1930 236 1933 303
rect 1922 233 1933 236
rect 1946 236 1949 323
rect 1946 233 1957 236
rect 1922 213 1925 233
rect 1866 203 1885 206
rect 1866 123 1869 203
rect 1914 193 1917 206
rect 1882 133 1885 146
rect 1930 123 1933 206
rect 1938 173 1941 216
rect 1946 183 1949 206
rect 1954 193 1957 233
rect 1962 213 1965 393
rect 1986 323 1989 513
rect 2018 476 2021 606
rect 2014 473 2021 476
rect 1994 413 1997 436
rect 2014 406 2017 473
rect 2026 413 2029 746
rect 2034 733 2037 816
rect 2042 783 2045 846
rect 2050 763 2053 906
rect 2058 756 2061 966
rect 2074 956 2077 1363
rect 2082 1323 2085 1406
rect 2082 963 2085 1316
rect 2090 1303 2093 1326
rect 2098 1323 2101 1426
rect 2114 1413 2117 1436
rect 2106 1393 2109 1406
rect 2106 1333 2109 1346
rect 2114 1233 2117 1406
rect 2122 1403 2125 1416
rect 2130 1413 2133 1426
rect 2122 1323 2125 1336
rect 2130 1306 2133 1406
rect 2138 1373 2141 1426
rect 2170 1383 2173 1726
rect 2194 1686 2197 1726
rect 2210 1706 2213 1806
rect 2246 1796 2249 1913
rect 2262 1906 2265 1973
rect 2242 1793 2249 1796
rect 2258 1903 2265 1906
rect 2242 1736 2245 1793
rect 2242 1733 2253 1736
rect 2250 1713 2253 1733
rect 2258 1723 2261 1903
rect 2210 1703 2217 1706
rect 2186 1683 2197 1686
rect 2178 1603 2181 1616
rect 2186 1603 2189 1683
rect 2214 1646 2217 1703
rect 2226 1656 2229 1676
rect 2226 1653 2233 1656
rect 2214 1643 2221 1646
rect 2202 1603 2205 1636
rect 2210 1613 2213 1626
rect 2186 1513 2189 1586
rect 2218 1563 2221 1643
rect 2230 1576 2233 1653
rect 2274 1623 2277 1976
rect 2282 1923 2285 1983
rect 2282 1716 2285 1886
rect 2290 1813 2293 1936
rect 2298 1883 2301 1956
rect 2306 1813 2309 1966
rect 2314 1933 2317 1946
rect 2322 1936 2325 2006
rect 2338 1993 2341 2006
rect 2338 1956 2341 1976
rect 2346 1963 2349 2016
rect 2354 2003 2357 2026
rect 2370 1973 2373 2156
rect 2378 2133 2381 2216
rect 2386 2193 2389 2233
rect 2386 2103 2389 2146
rect 2398 2096 2401 2243
rect 2410 2103 2413 2116
rect 2394 2093 2401 2096
rect 2394 2046 2397 2093
rect 2418 2086 2421 2353
rect 2426 2323 2429 2436
rect 2438 2426 2441 2483
rect 2450 2443 2453 2563
rect 2434 2423 2441 2426
rect 2434 2403 2437 2423
rect 2450 2413 2453 2426
rect 2458 2403 2461 2536
rect 2466 2433 2469 2716
rect 2482 2703 2485 2736
rect 2490 2713 2493 2736
rect 2474 2613 2477 2636
rect 2482 2526 2485 2606
rect 2490 2533 2493 2656
rect 2506 2603 2509 2746
rect 2530 2723 2533 2753
rect 2538 2733 2541 2816
rect 2546 2746 2549 2816
rect 2570 2813 2589 2816
rect 2554 2763 2557 2806
rect 2578 2803 2589 2806
rect 2594 2756 2597 2816
rect 2602 2813 2605 2823
rect 2578 2753 2597 2756
rect 2546 2743 2553 2746
rect 2538 2706 2541 2726
rect 2534 2703 2541 2706
rect 2534 2636 2537 2703
rect 2550 2696 2553 2743
rect 2578 2736 2581 2753
rect 2602 2746 2605 2806
rect 2626 2803 2629 2853
rect 2634 2813 2637 2826
rect 2634 2793 2637 2806
rect 2546 2693 2553 2696
rect 2574 2733 2581 2736
rect 2586 2743 2605 2746
rect 2534 2633 2541 2636
rect 2538 2613 2541 2633
rect 2514 2533 2517 2556
rect 2482 2523 2501 2526
rect 2474 2426 2477 2486
rect 2466 2423 2477 2426
rect 2410 2083 2421 2086
rect 2394 2043 2401 2046
rect 2398 1986 2401 2043
rect 2398 1983 2405 1986
rect 2338 1953 2349 1956
rect 2322 1933 2333 1936
rect 2346 1933 2349 1953
rect 2322 1913 2325 1926
rect 2370 1923 2373 1946
rect 2322 1813 2325 1826
rect 2338 1816 2341 1836
rect 2330 1813 2341 1816
rect 2346 1813 2365 1816
rect 2370 1813 2373 1836
rect 2298 1803 2309 1806
rect 2298 1753 2301 1803
rect 2314 1793 2317 1806
rect 2330 1803 2341 1806
rect 2282 1713 2293 1716
rect 2290 1666 2293 1713
rect 2286 1663 2293 1666
rect 2286 1616 2289 1663
rect 2230 1573 2237 1576
rect 2250 1573 2253 1616
rect 2282 1613 2289 1616
rect 2298 1613 2301 1626
rect 2194 1513 2197 1536
rect 2210 1533 2213 1556
rect 2218 1533 2221 1546
rect 2234 1526 2237 1573
rect 2282 1556 2285 1613
rect 2314 1603 2317 1726
rect 2322 1623 2325 1736
rect 2250 1533 2253 1546
rect 2202 1506 2205 1526
rect 2210 1513 2213 1526
rect 2226 1523 2237 1526
rect 2194 1503 2205 1506
rect 2194 1423 2197 1503
rect 2202 1413 2205 1496
rect 2126 1303 2133 1306
rect 2090 1213 2093 1226
rect 2126 1216 2129 1303
rect 2126 1213 2133 1216
rect 2130 1193 2133 1213
rect 2098 1133 2101 1156
rect 2090 1106 2093 1126
rect 2090 1103 2097 1106
rect 2094 1036 2097 1103
rect 2106 1063 2109 1176
rect 2138 1173 2141 1366
rect 2194 1346 2197 1406
rect 2210 1393 2213 1486
rect 2194 1343 2205 1346
rect 2146 1223 2149 1336
rect 2154 1213 2157 1326
rect 2162 1303 2165 1326
rect 2178 1286 2181 1336
rect 2202 1323 2205 1343
rect 2178 1283 2189 1286
rect 2170 1223 2173 1236
rect 2146 1156 2149 1206
rect 2138 1153 2149 1156
rect 2114 1133 2117 1146
rect 2122 1106 2125 1126
rect 2118 1103 2125 1106
rect 2090 1033 2097 1036
rect 2118 1036 2121 1103
rect 2118 1033 2125 1036
rect 2090 1013 2093 1033
rect 2122 1013 2125 1033
rect 2098 986 2101 1006
rect 2094 983 2101 986
rect 2066 953 2077 956
rect 2066 893 2069 953
rect 2074 923 2077 946
rect 2094 916 2097 983
rect 2122 976 2125 1006
rect 2106 973 2125 976
rect 2106 923 2109 973
rect 2094 913 2101 916
rect 2074 803 2077 856
rect 2034 523 2037 566
rect 2034 413 2037 426
rect 2014 403 2021 406
rect 2018 333 2021 403
rect 2034 343 2037 406
rect 2042 403 2045 756
rect 2050 753 2061 756
rect 2050 696 2053 753
rect 2082 743 2085 816
rect 2066 713 2069 736
rect 2050 693 2057 696
rect 2054 636 2057 693
rect 2050 633 2057 636
rect 2050 453 2053 633
rect 2058 606 2061 616
rect 2066 613 2069 636
rect 2058 603 2069 606
rect 2066 583 2069 603
rect 2058 433 2061 536
rect 2074 516 2077 686
rect 2082 623 2085 646
rect 2090 613 2093 826
rect 2098 793 2101 913
rect 2114 906 2117 956
rect 2110 903 2117 906
rect 2110 826 2113 903
rect 2106 823 2113 826
rect 2090 586 2093 606
rect 2098 603 2101 776
rect 2106 706 2109 823
rect 2114 773 2117 816
rect 2122 813 2125 966
rect 2130 953 2133 1136
rect 2138 1113 2141 1153
rect 2130 933 2133 946
rect 2130 916 2133 926
rect 2138 923 2141 1016
rect 2146 1013 2149 1026
rect 2154 1003 2157 1206
rect 2170 1193 2173 1206
rect 2186 1186 2189 1283
rect 2210 1193 2213 1216
rect 2178 1183 2189 1186
rect 2162 1133 2165 1146
rect 2178 1133 2181 1183
rect 2218 1176 2221 1386
rect 2226 1353 2229 1523
rect 2250 1256 2253 1526
rect 2258 1323 2261 1556
rect 2266 1553 2285 1556
rect 2266 1403 2269 1553
rect 2274 1513 2277 1536
rect 2290 1533 2293 1566
rect 2314 1523 2317 1546
rect 2330 1536 2333 1746
rect 2338 1633 2341 1736
rect 2346 1613 2349 1806
rect 2354 1733 2357 1806
rect 2354 1566 2357 1726
rect 2362 1716 2365 1813
rect 2370 1733 2373 1806
rect 2386 1783 2389 1976
rect 2402 1973 2405 1983
rect 2410 1923 2413 2083
rect 2426 2056 2429 2256
rect 2434 2133 2437 2326
rect 2458 2323 2461 2396
rect 2458 2253 2461 2316
rect 2466 2246 2469 2336
rect 2474 2303 2477 2423
rect 2482 2333 2485 2406
rect 2490 2316 2493 2446
rect 2498 2396 2501 2426
rect 2514 2413 2517 2526
rect 2538 2416 2541 2526
rect 2546 2523 2549 2693
rect 2554 2566 2557 2646
rect 2574 2596 2577 2733
rect 2586 2683 2589 2743
rect 2594 2676 2597 2736
rect 2610 2733 2621 2736
rect 2602 2713 2605 2726
rect 2626 2723 2629 2786
rect 2650 2783 2653 2816
rect 2658 2803 2661 2826
rect 2690 2823 2693 2856
rect 2698 2836 2701 2926
rect 2762 2853 2765 2926
rect 2778 2923 2781 2936
rect 2698 2833 2709 2836
rect 2770 2833 2773 2916
rect 2818 2866 2821 3040
rect 2858 2933 2861 2946
rect 2810 2863 2821 2866
rect 2634 2733 2637 2746
rect 2586 2673 2597 2676
rect 2586 2606 2589 2673
rect 2594 2613 2597 2626
rect 2586 2603 2597 2606
rect 2574 2593 2581 2596
rect 2554 2563 2561 2566
rect 2558 2516 2561 2563
rect 2554 2513 2561 2516
rect 2530 2413 2541 2416
rect 2546 2413 2549 2426
rect 2522 2396 2525 2406
rect 2530 2403 2533 2413
rect 2498 2393 2509 2396
rect 2522 2393 2533 2396
rect 2554 2393 2557 2513
rect 2562 2423 2565 2456
rect 2506 2346 2509 2393
rect 2498 2343 2509 2346
rect 2498 2323 2501 2343
rect 2530 2336 2533 2393
rect 2522 2333 2533 2336
rect 2482 2293 2485 2316
rect 2490 2313 2501 2316
rect 2498 2256 2501 2313
rect 2522 2266 2525 2333
rect 2522 2263 2533 2266
rect 2494 2253 2501 2256
rect 2466 2243 2477 2246
rect 2450 2203 2453 2216
rect 2426 2053 2445 2056
rect 2418 1993 2421 2016
rect 2426 1906 2429 1956
rect 2418 1903 2429 1906
rect 2418 1836 2421 1903
rect 2418 1833 2425 1836
rect 2410 1793 2413 1816
rect 2362 1713 2369 1716
rect 2366 1646 2369 1713
rect 2386 1686 2389 1766
rect 2410 1723 2413 1736
rect 2422 1706 2425 1833
rect 2422 1703 2429 1706
rect 2386 1683 2405 1686
rect 2426 1683 2429 1703
rect 2362 1643 2369 1646
rect 2362 1603 2365 1643
rect 2370 1603 2373 1626
rect 2378 1613 2381 1636
rect 2386 1603 2389 1616
rect 2354 1563 2361 1566
rect 2326 1533 2333 1536
rect 2314 1423 2317 1436
rect 2274 1383 2277 1416
rect 2306 1393 2309 1416
rect 2314 1383 2317 1406
rect 2326 1396 2329 1533
rect 2326 1393 2333 1396
rect 2274 1303 2277 1326
rect 2250 1253 2261 1256
rect 2214 1173 2221 1176
rect 2202 1123 2205 1146
rect 2162 1103 2165 1116
rect 2178 1066 2181 1116
rect 2214 1076 2217 1173
rect 2226 1083 2229 1246
rect 2258 1176 2261 1253
rect 2274 1223 2277 1296
rect 2282 1283 2285 1376
rect 2330 1373 2333 1393
rect 2298 1333 2301 1356
rect 2274 1206 2277 1216
rect 2282 1213 2285 1236
rect 2314 1223 2317 1286
rect 2274 1203 2293 1206
rect 2250 1173 2261 1176
rect 2250 1093 2253 1173
rect 2258 1133 2269 1136
rect 2290 1133 2293 1203
rect 2298 1183 2301 1206
rect 2258 1113 2261 1133
rect 2266 1103 2269 1126
rect 2282 1096 2285 1116
rect 2298 1103 2301 1126
rect 2306 1123 2309 1216
rect 2314 1196 2317 1216
rect 2322 1203 2325 1326
rect 2314 1193 2325 1196
rect 2282 1093 2293 1096
rect 2306 1093 2309 1116
rect 2214 1073 2221 1076
rect 2178 1063 2185 1066
rect 2130 913 2137 916
rect 2134 836 2137 913
rect 2134 833 2141 836
rect 2122 766 2125 806
rect 2130 803 2133 816
rect 2138 783 2141 833
rect 2146 813 2149 956
rect 2154 903 2157 936
rect 2146 793 2149 806
rect 2114 763 2125 766
rect 2114 723 2117 763
rect 2106 703 2117 706
rect 2106 593 2109 606
rect 2114 586 2117 703
rect 2122 613 2125 626
rect 2090 583 2117 586
rect 2070 513 2077 516
rect 2070 436 2073 513
rect 2070 433 2077 436
rect 2050 413 2061 416
rect 1970 203 1981 206
rect 1986 183 1989 216
rect 1994 213 1997 226
rect 2010 183 2013 326
rect 2034 323 2037 336
rect 2034 203 2037 216
rect 2050 213 2053 346
rect 2058 333 2061 406
rect 2066 326 2069 416
rect 2074 343 2077 433
rect 2082 423 2085 536
rect 2098 533 2101 583
rect 2122 566 2125 606
rect 2138 576 2141 716
rect 2154 706 2157 896
rect 2162 843 2165 1006
rect 2170 853 2173 1056
rect 2182 966 2185 1063
rect 2218 1053 2221 1073
rect 2282 1066 2285 1086
rect 2278 1063 2285 1066
rect 2290 1066 2293 1093
rect 2290 1063 2301 1066
rect 2194 1023 2197 1036
rect 2194 993 2197 1006
rect 2178 963 2185 966
rect 2178 926 2181 963
rect 2210 956 2213 1006
rect 2234 993 2237 1016
rect 2278 976 2281 1063
rect 2298 1026 2301 1063
rect 2290 1023 2301 1026
rect 2278 973 2285 976
rect 2210 953 2221 956
rect 2186 933 2189 946
rect 2178 923 2189 926
rect 2202 923 2205 936
rect 2186 826 2189 923
rect 2186 823 2213 826
rect 2162 733 2165 806
rect 2170 713 2173 806
rect 2178 783 2181 806
rect 2186 723 2189 806
rect 2194 716 2197 816
rect 2202 783 2205 806
rect 2210 766 2213 823
rect 2218 813 2221 953
rect 2242 923 2245 946
rect 2226 823 2229 886
rect 2226 793 2229 806
rect 2242 803 2245 816
rect 2266 793 2269 816
rect 2186 713 2197 716
rect 2202 763 2213 766
rect 2154 703 2173 706
rect 2170 636 2173 703
rect 2170 633 2177 636
rect 2162 593 2165 616
rect 2130 566 2133 576
rect 2138 573 2149 576
rect 2122 563 2133 566
rect 2090 473 2093 526
rect 2106 443 2109 536
rect 2114 533 2117 546
rect 2130 533 2133 563
rect 2130 513 2133 526
rect 2146 523 2149 573
rect 2174 566 2177 633
rect 2186 573 2189 713
rect 2202 643 2205 763
rect 2242 746 2245 786
rect 2234 743 2245 746
rect 2218 723 2221 736
rect 2234 696 2237 743
rect 2234 693 2245 696
rect 2234 613 2237 626
rect 2174 563 2181 566
rect 2170 523 2173 546
rect 2178 533 2181 563
rect 2242 536 2245 693
rect 2266 676 2269 736
rect 2282 733 2285 973
rect 2290 936 2293 1023
rect 2298 1006 2301 1016
rect 2306 1013 2309 1036
rect 2314 1006 2317 1136
rect 2322 1123 2325 1193
rect 2298 1003 2317 1006
rect 2322 1003 2325 1116
rect 2330 1096 2333 1236
rect 2338 1213 2341 1526
rect 2358 1486 2361 1563
rect 2370 1513 2373 1586
rect 2402 1573 2405 1683
rect 2426 1613 2429 1626
rect 2434 1583 2437 2026
rect 2442 1996 2445 2053
rect 2450 2013 2453 2196
rect 2458 2133 2461 2176
rect 2458 2023 2461 2126
rect 2442 1993 2453 1996
rect 2458 1993 2461 2006
rect 2450 1986 2453 1993
rect 2442 1976 2445 1986
rect 2450 1983 2461 1986
rect 2442 1973 2453 1976
rect 2442 1913 2445 1946
rect 2450 1933 2453 1973
rect 2450 1726 2453 1926
rect 2458 1743 2461 1983
rect 2466 1823 2469 2126
rect 2474 2116 2477 2243
rect 2482 2133 2485 2216
rect 2494 2196 2497 2253
rect 2494 2193 2501 2196
rect 2490 2133 2493 2176
rect 2498 2126 2501 2193
rect 2514 2176 2517 2236
rect 2490 2123 2501 2126
rect 2506 2173 2517 2176
rect 2530 2173 2533 2263
rect 2538 2223 2541 2236
rect 2474 2113 2481 2116
rect 2478 2046 2481 2113
rect 2474 2043 2481 2046
rect 2474 2023 2477 2043
rect 2474 1943 2477 2016
rect 2482 1936 2485 2006
rect 2490 1983 2493 2123
rect 2498 2013 2501 2026
rect 2506 2023 2509 2173
rect 2538 2166 2541 2216
rect 2514 2133 2517 2146
rect 2474 1933 2485 1936
rect 2498 1933 2501 2006
rect 2450 1723 2457 1726
rect 2466 1723 2469 1736
rect 2378 1523 2381 1536
rect 2402 1523 2405 1536
rect 2378 1513 2389 1516
rect 2354 1483 2361 1486
rect 2346 1393 2349 1406
rect 2354 1363 2357 1483
rect 2346 1213 2349 1256
rect 2354 1213 2357 1266
rect 2362 1213 2365 1236
rect 2370 1166 2373 1496
rect 2410 1446 2413 1556
rect 2426 1533 2429 1546
rect 2434 1533 2437 1556
rect 2402 1443 2413 1446
rect 2394 1383 2397 1416
rect 2402 1403 2405 1443
rect 2402 1333 2405 1356
rect 2394 1253 2397 1326
rect 2410 1323 2413 1416
rect 2418 1326 2421 1436
rect 2434 1413 2437 1526
rect 2442 1493 2445 1686
rect 2454 1666 2457 1723
rect 2474 1706 2477 1926
rect 2482 1846 2485 1933
rect 2498 1916 2501 1926
rect 2506 1923 2509 2016
rect 2498 1913 2509 1916
rect 2482 1843 2509 1846
rect 2482 1813 2485 1826
rect 2490 1813 2493 1836
rect 2506 1813 2509 1843
rect 2514 1833 2517 2126
rect 2522 2106 2525 2166
rect 2530 2163 2541 2166
rect 2546 2163 2549 2326
rect 2530 2126 2533 2163
rect 2554 2153 2557 2336
rect 2562 2213 2565 2416
rect 2570 2393 2573 2406
rect 2578 2396 2581 2593
rect 2586 2403 2589 2536
rect 2594 2403 2597 2596
rect 2602 2513 2605 2666
rect 2610 2643 2613 2716
rect 2650 2703 2653 2776
rect 2666 2763 2669 2806
rect 2674 2743 2677 2816
rect 2690 2803 2693 2816
rect 2706 2813 2709 2833
rect 2706 2773 2709 2806
rect 2730 2803 2733 2816
rect 2802 2813 2805 2826
rect 2794 2766 2797 2806
rect 2810 2803 2813 2863
rect 2826 2813 2829 2836
rect 2834 2803 2837 2926
rect 2858 2816 2861 2926
rect 2874 2836 2877 2926
rect 2882 2923 2885 2936
rect 2914 2933 2917 2946
rect 2930 2933 2933 2956
rect 2954 2923 2957 2946
rect 2866 2833 2877 2836
rect 2866 2823 2869 2833
rect 2786 2763 2797 2766
rect 2674 2723 2677 2736
rect 2610 2566 2613 2616
rect 2626 2613 2629 2636
rect 2634 2613 2637 2626
rect 2618 2593 2621 2606
rect 2642 2603 2645 2686
rect 2610 2563 2621 2566
rect 2578 2393 2589 2396
rect 2602 2393 2605 2416
rect 2570 2323 2573 2376
rect 2570 2293 2573 2316
rect 2578 2213 2581 2336
rect 2586 2213 2589 2393
rect 2594 2323 2597 2386
rect 2562 2193 2565 2206
rect 2594 2166 2597 2316
rect 2610 2233 2613 2556
rect 2618 2533 2621 2563
rect 2618 2496 2621 2526
rect 2626 2513 2629 2546
rect 2650 2533 2653 2616
rect 2634 2506 2637 2526
rect 2658 2523 2661 2626
rect 2666 2613 2669 2636
rect 2674 2613 2677 2626
rect 2674 2593 2677 2606
rect 2682 2603 2685 2616
rect 2682 2533 2685 2576
rect 2690 2533 2693 2616
rect 2690 2506 2693 2526
rect 2634 2503 2645 2506
rect 2618 2493 2625 2496
rect 2622 2366 2625 2493
rect 2642 2436 2645 2503
rect 2682 2503 2693 2506
rect 2634 2433 2645 2436
rect 2634 2403 2637 2433
rect 2622 2363 2637 2366
rect 2634 2313 2637 2363
rect 2586 2163 2597 2166
rect 2538 2133 2541 2146
rect 2530 2123 2541 2126
rect 2538 2113 2541 2123
rect 2522 2103 2529 2106
rect 2526 2036 2529 2103
rect 2554 2076 2557 2136
rect 2578 2123 2581 2146
rect 2554 2073 2565 2076
rect 2522 2033 2529 2036
rect 2522 1883 2525 2033
rect 2530 1933 2533 2016
rect 2538 1953 2541 2026
rect 2546 1993 2549 2006
rect 2562 1986 2565 2073
rect 2586 2023 2589 2163
rect 2586 2003 2589 2016
rect 2594 1993 2597 2156
rect 2554 1983 2565 1986
rect 2538 1933 2541 1946
rect 2530 1823 2533 1926
rect 2538 1896 2541 1916
rect 2538 1893 2545 1896
rect 2542 1826 2545 1893
rect 2538 1823 2545 1826
rect 2450 1663 2457 1666
rect 2470 1703 2477 1706
rect 2450 1576 2453 1663
rect 2470 1636 2473 1703
rect 2470 1633 2477 1636
rect 2474 1613 2477 1633
rect 2482 1613 2485 1736
rect 2490 1733 2493 1806
rect 2514 1803 2517 1816
rect 2538 1803 2541 1823
rect 2546 1786 2549 1806
rect 2538 1783 2549 1786
rect 2490 1696 2493 1716
rect 2490 1693 2497 1696
rect 2494 1626 2497 1693
rect 2506 1683 2509 1736
rect 2538 1716 2541 1783
rect 2554 1763 2557 1983
rect 2602 1966 2605 2216
rect 2618 2123 2621 2216
rect 2626 2116 2629 2206
rect 2634 2123 2637 2226
rect 2642 2213 2645 2416
rect 2650 2413 2661 2416
rect 2666 2413 2669 2466
rect 2682 2446 2685 2503
rect 2682 2443 2693 2446
rect 2674 2413 2677 2426
rect 2690 2413 2693 2443
rect 2626 2113 2637 2116
rect 2610 2003 2613 2066
rect 2626 1966 2629 2106
rect 2594 1963 2605 1966
rect 2622 1963 2629 1966
rect 2578 1913 2581 1926
rect 2594 1886 2597 1963
rect 2622 1916 2625 1963
rect 2634 1923 2637 2113
rect 2642 2106 2645 2206
rect 2650 2203 2653 2406
rect 2658 2366 2661 2413
rect 2698 2406 2701 2606
rect 2706 2523 2709 2636
rect 2714 2613 2717 2746
rect 2730 2656 2733 2726
rect 2722 2653 2733 2656
rect 2722 2573 2725 2653
rect 2714 2523 2717 2536
rect 2722 2533 2725 2546
rect 2730 2516 2733 2626
rect 2690 2403 2701 2406
rect 2658 2363 2677 2366
rect 2658 2323 2661 2346
rect 2658 2193 2661 2316
rect 2674 2306 2677 2363
rect 2690 2323 2693 2403
rect 2706 2343 2709 2406
rect 2714 2373 2717 2516
rect 2726 2513 2733 2516
rect 2726 2426 2729 2513
rect 2722 2423 2729 2426
rect 2738 2423 2741 2606
rect 2746 2553 2749 2736
rect 2770 2616 2773 2726
rect 2786 2686 2789 2763
rect 2834 2736 2837 2766
rect 2834 2733 2845 2736
rect 2786 2683 2797 2686
rect 2762 2613 2773 2616
rect 2762 2603 2765 2613
rect 2778 2603 2781 2616
rect 2794 2613 2797 2683
rect 2826 2676 2829 2726
rect 2834 2693 2837 2726
rect 2818 2673 2829 2676
rect 2818 2616 2821 2673
rect 2818 2613 2829 2616
rect 2794 2593 2797 2606
rect 2826 2593 2829 2613
rect 2842 2606 2845 2733
rect 2850 2713 2853 2816
rect 2858 2813 2869 2816
rect 2858 2733 2861 2796
rect 2866 2733 2869 2813
rect 2858 2713 2861 2726
rect 2866 2653 2869 2726
rect 2874 2716 2877 2826
rect 2882 2723 2885 2816
rect 2890 2803 2893 2826
rect 2898 2813 2901 2826
rect 2906 2806 2909 2866
rect 2914 2813 2917 2916
rect 3010 2863 3013 2926
rect 2906 2803 2917 2806
rect 2898 2733 2901 2746
rect 2874 2713 2901 2716
rect 2914 2713 2917 2736
rect 2898 2626 2901 2713
rect 2874 2623 2901 2626
rect 2842 2603 2869 2606
rect 2746 2503 2749 2536
rect 2762 2533 2765 2556
rect 2786 2523 2789 2546
rect 2842 2533 2853 2536
rect 2842 2526 2845 2533
rect 2834 2523 2845 2526
rect 2850 2503 2853 2526
rect 2834 2423 2853 2426
rect 2722 2383 2725 2423
rect 2730 2403 2733 2416
rect 2738 2343 2741 2416
rect 2746 2363 2749 2406
rect 2778 2393 2781 2416
rect 2802 2393 2805 2406
rect 2706 2323 2709 2336
rect 2674 2303 2685 2306
rect 2666 2203 2669 2266
rect 2682 2236 2685 2303
rect 2674 2233 2685 2236
rect 2674 2213 2677 2233
rect 2682 2213 2693 2216
rect 2666 2193 2685 2196
rect 2650 2123 2653 2136
rect 2658 2133 2661 2146
rect 2642 2103 2649 2106
rect 2646 2026 2649 2103
rect 2646 2023 2653 2026
rect 2642 1993 2645 2016
rect 2650 2003 2653 2023
rect 2658 1976 2661 2126
rect 2666 2046 2669 2126
rect 2674 2066 2677 2136
rect 2682 2133 2685 2193
rect 2690 2126 2693 2206
rect 2698 2203 2701 2306
rect 2730 2303 2733 2326
rect 2706 2223 2709 2246
rect 2706 2153 2709 2216
rect 2682 2123 2693 2126
rect 2698 2123 2701 2136
rect 2674 2063 2685 2066
rect 2666 2043 2673 2046
rect 2650 1973 2661 1976
rect 2650 1926 2653 1973
rect 2670 1956 2673 2043
rect 2682 2003 2685 2063
rect 2666 1953 2673 1956
rect 2666 1933 2669 1953
rect 2650 1923 2661 1926
rect 2622 1913 2629 1916
rect 2562 1813 2565 1886
rect 2594 1883 2605 1886
rect 2554 1723 2557 1746
rect 2538 1713 2549 1716
rect 2546 1686 2549 1713
rect 2538 1683 2549 1686
rect 2538 1636 2541 1683
rect 2538 1633 2549 1636
rect 2490 1623 2497 1626
rect 2490 1593 2493 1623
rect 2450 1573 2461 1576
rect 2450 1533 2453 1546
rect 2450 1473 2453 1526
rect 2458 1423 2461 1573
rect 2498 1553 2501 1606
rect 2426 1393 2429 1406
rect 2426 1333 2429 1376
rect 2450 1346 2453 1406
rect 2458 1403 2461 1416
rect 2482 1406 2485 1526
rect 2498 1523 2501 1546
rect 2506 1516 2509 1606
rect 2514 1603 2517 1616
rect 2546 1536 2549 1633
rect 2562 1596 2565 1686
rect 2578 1603 2581 1816
rect 2602 1803 2605 1883
rect 2618 1813 2621 1836
rect 2626 1806 2629 1913
rect 2658 1816 2661 1923
rect 2674 1913 2677 1926
rect 2682 1853 2685 1936
rect 2690 1846 2693 2036
rect 2698 1933 2701 2086
rect 2706 2013 2709 2136
rect 2714 2133 2717 2206
rect 2722 2203 2725 2216
rect 2738 2203 2741 2236
rect 2714 2106 2717 2126
rect 2722 2123 2725 2196
rect 2714 2103 2721 2106
rect 2730 2103 2733 2156
rect 2738 2133 2741 2146
rect 2778 2133 2781 2216
rect 2786 2153 2789 2326
rect 2802 2323 2805 2336
rect 2826 2323 2829 2406
rect 2866 2393 2869 2603
rect 2874 2593 2877 2606
rect 2890 2526 2893 2623
rect 2914 2603 2917 2616
rect 2898 2533 2901 2546
rect 2890 2523 2901 2526
rect 2914 2523 2917 2536
rect 2898 2423 2901 2523
rect 2718 2026 2721 2103
rect 2714 2023 2721 2026
rect 2746 2023 2749 2046
rect 2714 1953 2717 2023
rect 2730 2013 2741 2016
rect 2706 1933 2709 1946
rect 2682 1843 2693 1846
rect 2618 1803 2629 1806
rect 2650 1813 2669 1816
rect 2594 1733 2597 1746
rect 2586 1713 2589 1726
rect 2586 1613 2589 1626
rect 2594 1616 2597 1716
rect 2610 1703 2613 1726
rect 2594 1613 2605 1616
rect 2562 1593 2581 1596
rect 2498 1513 2509 1516
rect 2538 1533 2549 1536
rect 2578 1533 2581 1593
rect 2490 1413 2493 1426
rect 2482 1403 2493 1406
rect 2490 1393 2493 1403
rect 2498 1386 2501 1513
rect 2434 1333 2437 1346
rect 2442 1343 2453 1346
rect 2490 1383 2501 1386
rect 2418 1323 2429 1326
rect 2426 1313 2429 1323
rect 2434 1303 2437 1316
rect 2442 1253 2445 1343
rect 2386 1193 2389 1206
rect 2370 1163 2381 1166
rect 2338 1123 2341 1146
rect 2330 1093 2341 1096
rect 2338 1023 2341 1093
rect 2378 1086 2381 1163
rect 2370 1083 2381 1086
rect 2346 1013 2349 1056
rect 2370 1046 2373 1083
rect 2370 1043 2381 1046
rect 2290 933 2309 936
rect 2290 923 2301 926
rect 2306 856 2309 933
rect 2314 883 2317 926
rect 2306 853 2313 856
rect 2310 776 2313 853
rect 2322 813 2325 936
rect 2338 923 2341 1006
rect 2362 996 2365 1036
rect 2354 993 2365 996
rect 2354 936 2357 993
rect 2378 986 2381 1043
rect 2394 1003 2397 1126
rect 2418 1013 2421 1196
rect 2434 1176 2437 1216
rect 2450 1183 2453 1336
rect 2458 1313 2461 1326
rect 2434 1173 2453 1176
rect 2434 1133 2437 1146
rect 2434 1003 2437 1126
rect 2442 1123 2445 1166
rect 2450 1133 2453 1173
rect 2450 1113 2453 1126
rect 2458 1106 2461 1256
rect 2466 1213 2469 1336
rect 2490 1333 2493 1383
rect 2506 1353 2509 1476
rect 2538 1446 2541 1533
rect 2538 1443 2549 1446
rect 2514 1423 2517 1436
rect 2514 1413 2533 1416
rect 2514 1363 2517 1406
rect 2538 1403 2541 1426
rect 2546 1413 2549 1443
rect 2554 1413 2557 1526
rect 2474 1246 2477 1326
rect 2514 1323 2517 1346
rect 2474 1243 2485 1246
rect 2474 1223 2477 1236
rect 2474 1193 2477 1206
rect 2482 1176 2485 1243
rect 2466 1173 2485 1176
rect 2466 1123 2469 1173
rect 2490 1136 2493 1256
rect 2522 1253 2525 1376
rect 2538 1346 2541 1366
rect 2534 1343 2541 1346
rect 2562 1343 2565 1486
rect 2602 1483 2605 1536
rect 2578 1413 2581 1446
rect 2534 1286 2537 1343
rect 2570 1336 2573 1406
rect 2578 1386 2581 1406
rect 2586 1393 2589 1416
rect 2594 1403 2597 1416
rect 2602 1413 2605 1426
rect 2610 1413 2613 1626
rect 2618 1533 2621 1803
rect 2634 1766 2637 1796
rect 2650 1786 2653 1813
rect 2626 1763 2637 1766
rect 2646 1783 2653 1786
rect 2626 1713 2629 1763
rect 2646 1716 2649 1783
rect 2658 1723 2661 1806
rect 2682 1766 2685 1843
rect 2690 1823 2693 1836
rect 2698 1813 2701 1926
rect 2714 1913 2717 1936
rect 2722 1923 2725 2006
rect 2738 1963 2741 2006
rect 2698 1793 2701 1806
rect 2682 1763 2693 1766
rect 2690 1746 2693 1763
rect 2690 1743 2697 1746
rect 2646 1713 2653 1716
rect 2626 1623 2629 1706
rect 2650 1696 2653 1713
rect 2650 1693 2661 1696
rect 2634 1613 2637 1626
rect 2618 1506 2621 1526
rect 2618 1503 2625 1506
rect 2622 1436 2625 1503
rect 2634 1473 2637 1526
rect 2642 1523 2645 1606
rect 2658 1603 2661 1693
rect 2694 1686 2697 1743
rect 2690 1683 2697 1686
rect 2666 1613 2669 1646
rect 2682 1606 2685 1626
rect 2678 1603 2685 1606
rect 2678 1446 2681 1603
rect 2690 1473 2693 1683
rect 2698 1613 2701 1636
rect 2698 1593 2701 1606
rect 2706 1553 2709 1856
rect 2714 1813 2717 1906
rect 2730 1803 2733 1946
rect 2738 1903 2741 1956
rect 2746 1923 2749 2006
rect 2754 2003 2757 2126
rect 2762 2113 2765 2126
rect 2762 2026 2765 2046
rect 2762 2023 2773 2026
rect 2778 2023 2781 2036
rect 2786 2026 2789 2136
rect 2802 2123 2805 2226
rect 2818 2136 2821 2216
rect 2834 2203 2837 2326
rect 2874 2303 2877 2416
rect 2882 2323 2885 2406
rect 2914 2403 2917 2426
rect 2890 2333 2893 2396
rect 2898 2323 2901 2346
rect 2914 2333 2917 2396
rect 2930 2323 2933 2806
rect 2954 2793 2957 2816
rect 3010 2813 3013 2826
rect 2954 2723 2957 2746
rect 3010 2713 3013 2736
rect 2954 2593 2957 2616
rect 3002 2613 3013 2616
rect 2954 2523 2957 2546
rect 3010 2526 3013 2536
rect 3002 2523 3013 2526
rect 2954 2393 2957 2416
rect 3010 2413 3013 2426
rect 2914 2303 2917 2316
rect 2810 2133 2821 2136
rect 2794 2113 2805 2116
rect 2794 2033 2797 2113
rect 2786 2023 2797 2026
rect 2762 2003 2765 2016
rect 2754 1873 2757 1986
rect 2762 1916 2765 1976
rect 2770 1923 2773 2023
rect 2778 1993 2781 2006
rect 2786 2003 2789 2016
rect 2786 1983 2789 1996
rect 2794 1993 2797 2023
rect 2762 1913 2773 1916
rect 2778 1913 2781 1926
rect 2738 1796 2741 1816
rect 2746 1813 2749 1826
rect 2762 1813 2765 1913
rect 2786 1886 2789 1956
rect 2770 1883 2789 1886
rect 2770 1813 2773 1883
rect 2778 1813 2781 1826
rect 2786 1806 2789 1876
rect 2794 1823 2797 1916
rect 2802 1816 2805 2096
rect 2810 2066 2813 2133
rect 2818 2083 2821 2126
rect 2826 2106 2829 2146
rect 2834 2126 2837 2196
rect 2858 2176 2861 2216
rect 2842 2173 2861 2176
rect 2842 2133 2845 2173
rect 2858 2133 2861 2166
rect 2834 2123 2845 2126
rect 2842 2113 2845 2123
rect 2826 2103 2833 2106
rect 2810 2063 2821 2066
rect 2810 1993 2813 2036
rect 2818 1966 2821 2063
rect 2830 2036 2833 2103
rect 2826 2033 2833 2036
rect 2826 2013 2829 2033
rect 2810 1963 2821 1966
rect 2810 1843 2813 1963
rect 2826 1953 2829 2006
rect 2826 1886 2829 1946
rect 2818 1883 2829 1886
rect 2794 1813 2805 1816
rect 2810 1813 2813 1826
rect 2786 1803 2797 1806
rect 2738 1793 2757 1796
rect 2714 1676 2717 1726
rect 2714 1673 2733 1676
rect 2698 1523 2701 1536
rect 2618 1433 2625 1436
rect 2674 1443 2681 1446
rect 2618 1413 2621 1433
rect 2626 1406 2629 1416
rect 2602 1403 2613 1406
rect 2618 1403 2629 1406
rect 2578 1383 2589 1386
rect 2558 1333 2573 1336
rect 2558 1286 2561 1333
rect 2534 1283 2541 1286
rect 2538 1226 2541 1283
rect 2554 1283 2561 1286
rect 2498 1213 2501 1226
rect 2538 1223 2549 1226
rect 2514 1173 2517 1206
rect 2538 1193 2541 1216
rect 2450 1103 2461 1106
rect 2450 1046 2453 1103
rect 2446 1043 2453 1046
rect 2370 983 2381 986
rect 2354 933 2365 936
rect 2362 916 2365 933
rect 2354 913 2365 916
rect 2330 803 2333 836
rect 2346 803 2349 866
rect 2354 783 2357 913
rect 2370 906 2373 983
rect 2446 936 2449 1043
rect 2474 1036 2477 1136
rect 2482 1126 2485 1136
rect 2490 1133 2501 1136
rect 2482 1123 2493 1126
rect 2482 1053 2485 1116
rect 2490 1096 2493 1123
rect 2498 1113 2501 1133
rect 2490 1093 2501 1096
rect 2458 1033 2477 1036
rect 2362 903 2373 906
rect 2362 823 2365 903
rect 2378 863 2381 916
rect 2370 813 2373 846
rect 2386 833 2389 936
rect 2446 933 2453 936
rect 2394 913 2397 926
rect 2410 923 2421 926
rect 2434 913 2445 916
rect 2450 896 2453 933
rect 2446 893 2453 896
rect 2378 823 2389 826
rect 2306 773 2313 776
rect 2282 713 2285 726
rect 2258 673 2269 676
rect 2258 576 2261 673
rect 2274 616 2277 686
rect 2306 683 2309 773
rect 2322 676 2325 736
rect 2330 683 2333 716
rect 2322 673 2333 676
rect 2274 613 2285 616
rect 2330 613 2333 673
rect 2362 653 2365 806
rect 2378 803 2381 816
rect 2370 716 2373 736
rect 2386 723 2389 816
rect 2426 813 2429 836
rect 2370 713 2377 716
rect 2394 713 2397 786
rect 2402 776 2405 806
rect 2402 773 2413 776
rect 2410 733 2413 773
rect 2434 746 2437 856
rect 2446 776 2449 893
rect 2458 853 2461 1033
rect 2474 943 2477 1016
rect 2498 1013 2501 1093
rect 2506 1023 2509 1136
rect 2514 1133 2517 1146
rect 2514 1103 2517 1116
rect 2530 1056 2533 1186
rect 2546 1153 2549 1223
rect 2538 1123 2541 1136
rect 2554 1133 2557 1283
rect 2570 1253 2573 1326
rect 2578 1226 2581 1376
rect 2586 1343 2589 1383
rect 2594 1333 2605 1336
rect 2610 1333 2613 1366
rect 2618 1333 2621 1403
rect 2586 1233 2589 1326
rect 2578 1223 2589 1226
rect 2586 1206 2589 1223
rect 2594 1213 2597 1226
rect 2602 1213 2605 1326
rect 2618 1293 2621 1316
rect 2626 1313 2629 1356
rect 2634 1323 2637 1336
rect 2650 1333 2653 1406
rect 2642 1306 2645 1326
rect 2638 1303 2645 1306
rect 2610 1213 2613 1236
rect 2618 1206 2621 1256
rect 2638 1236 2641 1303
rect 2638 1233 2645 1236
rect 2586 1203 2597 1206
rect 2610 1203 2621 1206
rect 2578 1123 2581 1146
rect 2586 1106 2589 1136
rect 2522 1053 2533 1056
rect 2582 1103 2589 1106
rect 2522 1036 2525 1053
rect 2518 1033 2525 1036
rect 2518 976 2521 1033
rect 2554 1006 2557 1016
rect 2562 1013 2565 1026
rect 2554 1003 2573 1006
rect 2570 993 2573 1003
rect 2582 986 2585 1103
rect 2582 983 2589 986
rect 2594 983 2597 1203
rect 2618 1173 2621 1203
rect 2602 1073 2605 1156
rect 2626 1143 2629 1226
rect 2634 1136 2637 1216
rect 2642 1213 2645 1233
rect 2650 1216 2653 1326
rect 2658 1323 2661 1356
rect 2666 1333 2669 1416
rect 2674 1333 2677 1443
rect 2698 1403 2701 1416
rect 2722 1413 2725 1616
rect 2730 1603 2733 1673
rect 2738 1613 2741 1736
rect 2754 1733 2757 1793
rect 2754 1636 2757 1656
rect 2770 1643 2773 1766
rect 2786 1733 2789 1746
rect 2794 1733 2797 1803
rect 2802 1783 2805 1813
rect 2818 1763 2821 1883
rect 2834 1846 2837 2016
rect 2842 2013 2845 2026
rect 2850 2006 2853 2126
rect 2866 2123 2869 2196
rect 2914 2186 2917 2216
rect 2922 2193 2925 2206
rect 2914 2183 2925 2186
rect 2914 2163 2917 2183
rect 2930 2156 2933 2216
rect 2954 2203 2957 2326
rect 2970 2166 2973 2236
rect 3010 2203 3013 2326
rect 2970 2163 2981 2166
rect 2930 2153 2941 2156
rect 2874 2123 2877 2146
rect 2890 2133 2893 2146
rect 2890 2103 2893 2116
rect 2866 2023 2869 2036
rect 2842 2003 2853 2006
rect 2842 1856 2845 1996
rect 2850 1973 2853 2003
rect 2866 1993 2869 2006
rect 2882 2003 2885 2056
rect 2906 2053 2909 2136
rect 2930 2123 2933 2146
rect 2938 2093 2941 2153
rect 2978 2116 2981 2163
rect 3010 2136 3013 2166
rect 2994 2133 3013 2136
rect 2994 2123 2997 2133
rect 2978 2113 2997 2116
rect 2930 2036 2933 2056
rect 2926 2033 2933 2036
rect 2850 1866 2853 1926
rect 2874 1903 2877 1936
rect 2890 1933 2893 1976
rect 2898 1923 2901 1966
rect 2850 1863 2869 1866
rect 2842 1853 2853 1856
rect 2834 1843 2845 1846
rect 2834 1816 2837 1826
rect 2826 1813 2837 1816
rect 2842 1813 2845 1843
rect 2810 1733 2813 1746
rect 2746 1633 2757 1636
rect 2754 1623 2757 1633
rect 2738 1593 2741 1606
rect 2738 1533 2741 1546
rect 2754 1443 2757 1566
rect 2762 1483 2765 1636
rect 2786 1633 2789 1716
rect 2786 1613 2789 1626
rect 2786 1593 2789 1606
rect 2794 1546 2797 1626
rect 2802 1613 2805 1646
rect 2810 1603 2813 1726
rect 2818 1546 2821 1626
rect 2826 1623 2829 1813
rect 2834 1793 2837 1806
rect 2842 1776 2845 1806
rect 2838 1773 2845 1776
rect 2838 1706 2841 1773
rect 2850 1716 2853 1853
rect 2858 1723 2861 1846
rect 2866 1813 2869 1863
rect 2906 1816 2909 2026
rect 2914 1993 2917 2016
rect 2926 1966 2929 2033
rect 2962 2006 2965 2016
rect 2970 2013 2973 2036
rect 2986 2023 2989 2113
rect 3002 2103 3005 2126
rect 2978 2006 2981 2016
rect 2962 2003 2981 2006
rect 2926 1963 2933 1966
rect 2914 1933 2917 1946
rect 2930 1933 2933 1963
rect 2914 1913 2917 1926
rect 2954 1923 2957 1946
rect 2994 1923 2997 2016
rect 3010 1923 3013 2006
rect 2914 1823 2917 1836
rect 2906 1813 2917 1816
rect 2874 1793 2877 1806
rect 2866 1723 2869 1746
rect 2874 1736 2877 1786
rect 2914 1746 2917 1813
rect 2898 1743 2917 1746
rect 2874 1733 2893 1736
rect 2874 1716 2877 1726
rect 2850 1713 2877 1716
rect 2838 1703 2845 1706
rect 2842 1643 2845 1703
rect 2770 1533 2781 1536
rect 2778 1513 2781 1526
rect 2730 1423 2749 1426
rect 2674 1313 2677 1326
rect 2666 1223 2669 1296
rect 2682 1293 2685 1346
rect 2690 1333 2693 1366
rect 2650 1213 2669 1216
rect 2618 1133 2637 1136
rect 2642 1133 2645 1206
rect 2618 1086 2621 1133
rect 2626 1123 2637 1126
rect 2610 1083 2621 1086
rect 2602 1013 2605 1026
rect 2610 1003 2613 1083
rect 2518 973 2525 976
rect 2474 926 2477 936
rect 2482 933 2493 936
rect 2498 926 2501 956
rect 2522 953 2525 973
rect 2586 966 2589 983
rect 2618 973 2621 1076
rect 2586 963 2593 966
rect 2466 913 2469 926
rect 2474 923 2485 926
rect 2490 923 2501 926
rect 2506 923 2509 936
rect 2482 813 2485 923
rect 2522 886 2525 946
rect 2546 923 2549 936
rect 2590 886 2593 963
rect 2522 883 2541 886
rect 2490 813 2493 826
rect 2514 813 2517 856
rect 2522 806 2525 826
rect 2446 773 2453 776
rect 2434 743 2441 746
rect 2374 616 2377 713
rect 2370 613 2377 616
rect 2386 613 2389 656
rect 2258 573 2269 576
rect 2274 573 2277 606
rect 2266 553 2269 573
rect 2282 556 2285 613
rect 2290 593 2293 606
rect 2274 553 2285 556
rect 2274 546 2277 553
rect 2266 543 2277 546
rect 2234 533 2245 536
rect 2106 423 2109 436
rect 2082 373 2085 406
rect 2090 403 2093 416
rect 2106 393 2109 406
rect 2106 333 2109 366
rect 2122 363 2125 406
rect 2146 393 2149 416
rect 2066 323 2085 326
rect 2154 323 2157 336
rect 2082 233 2085 323
rect 2106 213 2109 226
rect 2154 223 2165 226
rect 2170 213 2173 236
rect 2122 193 2125 206
rect 2130 203 2149 206
rect 1978 123 1981 176
rect 2082 133 2085 186
rect 2066 113 2069 126
rect 2130 123 2133 203
rect 2170 123 2173 206
rect 2178 193 2181 376
rect 2194 323 2197 346
rect 2202 333 2205 486
rect 2210 393 2213 416
rect 2218 413 2221 476
rect 2234 406 2237 533
rect 2242 513 2245 526
rect 2250 483 2253 536
rect 2266 526 2269 543
rect 2262 523 2269 526
rect 2274 523 2277 536
rect 2290 533 2293 556
rect 2306 553 2309 606
rect 2314 523 2317 576
rect 2262 446 2265 523
rect 2262 443 2269 446
rect 2266 413 2269 443
rect 2274 423 2277 516
rect 2282 413 2285 436
rect 2218 403 2237 406
rect 2234 376 2237 403
rect 2226 373 2237 376
rect 2226 326 2229 373
rect 2242 333 2245 406
rect 2250 343 2253 406
rect 2266 393 2269 406
rect 2202 313 2205 326
rect 2226 323 2237 326
rect 2234 233 2237 323
rect 2282 313 2285 336
rect 2226 223 2237 226
rect 2250 213 2253 246
rect 2282 206 2285 236
rect 2290 213 2293 426
rect 2306 413 2309 426
rect 2314 393 2317 406
rect 2314 333 2317 346
rect 2314 223 2317 236
rect 2322 213 2325 226
rect 2330 223 2333 556
rect 2354 413 2357 526
rect 2370 523 2373 613
rect 2394 583 2397 606
rect 2410 603 2413 726
rect 2438 696 2441 743
rect 2434 693 2441 696
rect 2434 636 2437 693
rect 2418 633 2437 636
rect 2418 613 2421 626
rect 2378 533 2381 566
rect 2394 526 2397 536
rect 2386 523 2397 526
rect 2386 453 2389 523
rect 2394 496 2397 516
rect 2402 503 2405 526
rect 2410 516 2413 586
rect 2418 523 2421 596
rect 2426 583 2429 633
rect 2434 623 2437 633
rect 2434 603 2437 616
rect 2442 613 2445 636
rect 2426 533 2429 546
rect 2442 523 2445 556
rect 2450 533 2453 773
rect 2458 723 2461 736
rect 2490 733 2493 806
rect 2506 803 2525 806
rect 2506 723 2509 803
rect 2514 733 2517 746
rect 2530 736 2533 826
rect 2538 753 2541 883
rect 2586 883 2593 886
rect 2546 813 2565 816
rect 2586 813 2589 883
rect 2602 863 2605 936
rect 2610 933 2613 956
rect 2626 933 2629 1046
rect 2642 1013 2645 1126
rect 2650 1123 2653 1136
rect 2658 1133 2661 1146
rect 2666 1036 2669 1213
rect 2650 1033 2669 1036
rect 2674 1033 2677 1216
rect 2682 1203 2685 1266
rect 2690 1203 2693 1326
rect 2698 1183 2701 1386
rect 2714 1353 2717 1406
rect 2706 1333 2709 1346
rect 2714 1303 2717 1336
rect 2722 1333 2725 1376
rect 2730 1333 2733 1416
rect 2738 1373 2741 1416
rect 2754 1393 2757 1426
rect 2762 1386 2765 1476
rect 2770 1393 2773 1406
rect 2778 1396 2781 1416
rect 2786 1403 2789 1546
rect 2794 1543 2805 1546
rect 2794 1513 2797 1536
rect 2802 1516 2805 1543
rect 2810 1543 2821 1546
rect 2810 1523 2813 1543
rect 2802 1513 2821 1516
rect 2778 1393 2789 1396
rect 2762 1383 2781 1386
rect 2730 1306 2733 1326
rect 2726 1303 2733 1306
rect 2650 1006 2653 1033
rect 2666 1023 2677 1026
rect 2610 923 2621 926
rect 2634 906 2637 1006
rect 2642 1003 2653 1006
rect 2642 916 2645 1003
rect 2658 996 2661 1016
rect 2666 1013 2677 1016
rect 2682 1013 2685 1126
rect 2690 1046 2693 1136
rect 2698 1133 2701 1176
rect 2698 1103 2701 1126
rect 2690 1043 2701 1046
rect 2706 1043 2709 1256
rect 2650 993 2661 996
rect 2650 933 2653 993
rect 2666 933 2669 986
rect 2674 933 2677 966
rect 2658 923 2677 926
rect 2642 913 2649 916
rect 2626 903 2637 906
rect 2626 836 2629 903
rect 2646 856 2649 913
rect 2674 906 2677 923
rect 2670 903 2677 906
rect 2646 853 2653 856
rect 2626 833 2637 836
rect 2546 803 2557 806
rect 2570 793 2573 806
rect 2522 733 2533 736
rect 2458 623 2461 646
rect 2482 613 2485 646
rect 2490 553 2493 656
rect 2506 623 2509 636
rect 2514 623 2517 716
rect 2522 686 2525 733
rect 2530 703 2533 726
rect 2538 713 2541 736
rect 2554 733 2557 756
rect 2578 723 2581 746
rect 2586 716 2589 806
rect 2610 803 2613 816
rect 2618 766 2621 816
rect 2618 763 2625 766
rect 2578 713 2589 716
rect 2522 683 2529 686
rect 2526 616 2529 683
rect 2578 626 2581 713
rect 2622 696 2625 763
rect 2618 693 2625 696
rect 2618 676 2621 693
rect 2610 673 2621 676
rect 2578 623 2589 626
rect 2522 613 2529 616
rect 2522 593 2525 613
rect 2538 596 2541 606
rect 2546 603 2557 606
rect 2538 593 2549 596
rect 2410 513 2421 516
rect 2410 496 2413 513
rect 2426 503 2429 516
rect 2394 493 2413 496
rect 2410 393 2413 456
rect 2442 406 2445 496
rect 2466 486 2469 536
rect 2490 523 2493 546
rect 2546 523 2549 593
rect 2554 533 2557 603
rect 2562 493 2565 616
rect 2586 576 2589 623
rect 2610 616 2613 673
rect 2634 656 2637 833
rect 2650 736 2653 853
rect 2658 776 2661 866
rect 2670 836 2673 903
rect 2670 833 2677 836
rect 2666 783 2669 816
rect 2674 793 2677 833
rect 2682 796 2685 1006
rect 2690 803 2693 1036
rect 2698 993 2701 1043
rect 2714 1033 2717 1216
rect 2726 1196 2729 1303
rect 2738 1253 2741 1366
rect 2746 1323 2749 1346
rect 2746 1303 2749 1316
rect 2738 1203 2741 1226
rect 2726 1193 2733 1196
rect 2722 1113 2725 1126
rect 2730 1116 2733 1193
rect 2746 1163 2749 1216
rect 2754 1213 2757 1336
rect 2770 1313 2773 1376
rect 2778 1333 2781 1383
rect 2778 1286 2781 1316
rect 2786 1303 2789 1393
rect 2770 1283 2781 1286
rect 2762 1213 2765 1226
rect 2754 1193 2757 1206
rect 2738 1143 2757 1146
rect 2738 1123 2741 1143
rect 2746 1123 2749 1136
rect 2754 1133 2757 1143
rect 2730 1113 2741 1116
rect 2706 1023 2733 1026
rect 2706 1013 2709 1023
rect 2698 813 2701 976
rect 2706 896 2709 966
rect 2714 933 2717 1016
rect 2722 1013 2733 1016
rect 2738 1013 2741 1113
rect 2754 1103 2757 1126
rect 2762 1033 2765 1206
rect 2770 1143 2773 1283
rect 2754 1023 2765 1026
rect 2770 1013 2773 1126
rect 2722 933 2725 1013
rect 2730 993 2733 1006
rect 2738 963 2741 1006
rect 2762 973 2765 1006
rect 2778 1003 2781 1276
rect 2786 1223 2789 1236
rect 2786 1133 2789 1216
rect 2794 1203 2797 1486
rect 2802 1313 2805 1506
rect 2818 1446 2821 1513
rect 2826 1506 2829 1616
rect 2834 1563 2837 1606
rect 2834 1533 2837 1546
rect 2842 1523 2845 1636
rect 2850 1623 2853 1636
rect 2858 1613 2861 1706
rect 2866 1623 2869 1713
rect 2874 1613 2877 1636
rect 2850 1593 2853 1606
rect 2882 1563 2885 1726
rect 2890 1613 2893 1733
rect 2898 1723 2901 1743
rect 2906 1733 2917 1736
rect 2898 1703 2901 1716
rect 2906 1693 2909 1726
rect 2914 1713 2917 1726
rect 2826 1503 2837 1506
rect 2814 1443 2821 1446
rect 2814 1356 2817 1443
rect 2834 1436 2837 1503
rect 2850 1493 2853 1556
rect 2866 1533 2869 1546
rect 2858 1523 2885 1526
rect 2866 1503 2869 1516
rect 2882 1473 2885 1523
rect 2890 1513 2893 1606
rect 2914 1603 2917 1626
rect 2930 1583 2933 1906
rect 3026 1883 3029 1916
rect 2946 1743 2949 1826
rect 2954 1723 2957 1806
rect 2954 1613 2957 1696
rect 2970 1656 2973 1736
rect 3010 1723 3013 1736
rect 2966 1653 2973 1656
rect 2930 1546 2933 1566
rect 2966 1556 2969 1653
rect 2978 1566 2981 1646
rect 2978 1563 2989 1566
rect 2966 1553 2973 1556
rect 2898 1496 2901 1546
rect 2926 1543 2933 1546
rect 2914 1513 2917 1526
rect 2826 1433 2837 1436
rect 2814 1353 2821 1356
rect 2810 1306 2813 1336
rect 2818 1323 2821 1353
rect 2802 1303 2813 1306
rect 2802 1203 2805 1303
rect 2810 1213 2813 1296
rect 2818 1213 2821 1316
rect 2794 1183 2797 1196
rect 2810 1146 2813 1206
rect 2818 1183 2821 1206
rect 2826 1146 2829 1433
rect 2834 1383 2837 1406
rect 2834 1333 2837 1366
rect 2834 1213 2837 1326
rect 2842 1206 2845 1416
rect 2850 1333 2853 1346
rect 2866 1333 2869 1406
rect 2874 1363 2877 1406
rect 2834 1203 2845 1206
rect 2850 1196 2853 1316
rect 2858 1306 2861 1326
rect 2858 1303 2865 1306
rect 2862 1226 2865 1303
rect 2846 1193 2853 1196
rect 2858 1223 2865 1226
rect 2802 1126 2805 1146
rect 2810 1143 2821 1146
rect 2826 1143 2837 1146
rect 2738 933 2741 946
rect 2754 933 2757 946
rect 2714 923 2725 926
rect 2714 913 2717 923
rect 2706 893 2717 896
rect 2714 826 2717 893
rect 2706 823 2717 826
rect 2730 823 2733 926
rect 2746 823 2749 836
rect 2682 793 2693 796
rect 2658 773 2669 776
rect 2642 733 2653 736
rect 2642 706 2645 733
rect 2650 713 2653 726
rect 2642 703 2653 706
rect 2634 653 2645 656
rect 2634 623 2637 646
rect 2610 613 2621 616
rect 2578 573 2589 576
rect 2578 523 2581 573
rect 2602 523 2605 536
rect 2618 513 2621 613
rect 2626 496 2629 526
rect 2466 483 2477 486
rect 2458 413 2461 436
rect 2418 383 2421 406
rect 2442 403 2461 406
rect 2474 403 2477 483
rect 2562 423 2565 436
rect 2354 313 2357 326
rect 2410 323 2413 346
rect 2418 333 2421 366
rect 2434 333 2437 346
rect 2434 313 2437 326
rect 2442 303 2445 326
rect 2458 313 2461 403
rect 2498 336 2501 416
rect 2482 333 2501 336
rect 2530 333 2533 376
rect 2554 373 2557 416
rect 2490 306 2493 326
rect 2482 303 2493 306
rect 2482 246 2485 303
rect 2498 293 2501 326
rect 2482 243 2493 246
rect 2194 133 2197 146
rect 2226 123 2229 206
rect 2274 123 2277 206
rect 2282 203 2293 206
rect 2290 133 2293 203
rect 2322 193 2325 206
rect 2330 166 2333 216
rect 2338 213 2341 236
rect 2346 213 2349 226
rect 2346 173 2349 206
rect 2362 183 2365 206
rect 2322 163 2333 166
rect 2282 113 2285 126
rect 2322 113 2325 163
rect 2330 133 2333 146
rect 2346 133 2349 156
rect 2378 153 2381 226
rect 2490 216 2493 243
rect 2402 193 2405 216
rect 2482 213 2493 216
rect 2498 213 2501 236
rect 2506 213 2509 246
rect 2514 213 2517 226
rect 2522 223 2525 236
rect 2530 223 2533 326
rect 2538 213 2541 296
rect 2546 286 2549 336
rect 2578 323 2581 406
rect 2594 366 2597 496
rect 2618 493 2629 496
rect 2618 426 2621 493
rect 2618 423 2629 426
rect 2590 363 2597 366
rect 2590 316 2593 363
rect 2626 323 2629 423
rect 2642 393 2645 653
rect 2650 533 2653 703
rect 2658 613 2661 726
rect 2666 623 2669 773
rect 2674 616 2677 756
rect 2666 613 2677 616
rect 2658 523 2661 606
rect 2666 506 2669 613
rect 2674 593 2677 606
rect 2682 546 2685 746
rect 2690 733 2693 793
rect 2698 783 2701 806
rect 2706 743 2709 823
rect 2730 813 2749 816
rect 2722 786 2725 806
rect 2722 783 2729 786
rect 2658 503 2669 506
rect 2674 543 2685 546
rect 2658 426 2661 503
rect 2658 423 2669 426
rect 2666 363 2669 423
rect 2674 383 2677 543
rect 2682 523 2685 536
rect 2682 403 2685 516
rect 2690 496 2693 636
rect 2698 613 2701 726
rect 2706 546 2709 736
rect 2714 733 2717 756
rect 2714 653 2717 726
rect 2726 706 2729 783
rect 2738 733 2741 806
rect 2746 796 2749 813
rect 2746 793 2757 796
rect 2746 723 2749 793
rect 2754 723 2757 736
rect 2762 733 2765 876
rect 2778 813 2781 926
rect 2786 806 2789 1036
rect 2794 1023 2797 1126
rect 2802 1123 2809 1126
rect 2806 1046 2809 1123
rect 2802 1043 2809 1046
rect 2802 1023 2805 1043
rect 2810 1006 2813 1016
rect 2794 1003 2813 1006
rect 2778 803 2789 806
rect 2778 733 2781 803
rect 2762 713 2765 726
rect 2786 723 2789 746
rect 2794 723 2797 986
rect 2802 876 2805 966
rect 2802 873 2809 876
rect 2806 816 2809 873
rect 2802 813 2809 816
rect 2802 733 2805 813
rect 2818 746 2821 1143
rect 2826 873 2829 1136
rect 2834 1093 2837 1143
rect 2846 1086 2849 1193
rect 2858 1133 2861 1223
rect 2858 1113 2861 1126
rect 2866 1086 2869 1206
rect 2874 1173 2877 1346
rect 2882 1213 2885 1386
rect 2890 1273 2893 1496
rect 2898 1493 2909 1496
rect 2906 1426 2909 1493
rect 2926 1446 2929 1543
rect 2926 1443 2933 1446
rect 2898 1423 2909 1426
rect 2898 1406 2901 1423
rect 2922 1413 2925 1426
rect 2898 1403 2925 1406
rect 2842 1083 2849 1086
rect 2858 1083 2869 1086
rect 2834 923 2837 1006
rect 2842 983 2845 1083
rect 2850 1013 2853 1026
rect 2842 916 2845 946
rect 2850 933 2853 1006
rect 2858 926 2861 1083
rect 2834 913 2845 916
rect 2850 923 2861 926
rect 2834 866 2837 913
rect 2810 743 2821 746
rect 2826 863 2837 866
rect 2726 703 2733 706
rect 2730 656 2733 703
rect 2810 693 2813 743
rect 2826 736 2829 863
rect 2834 773 2837 806
rect 2842 783 2845 806
rect 2818 733 2829 736
rect 2722 653 2733 656
rect 2722 633 2725 653
rect 2706 543 2717 546
rect 2698 513 2701 526
rect 2706 523 2709 536
rect 2714 516 2717 543
rect 2722 523 2725 626
rect 2706 513 2717 516
rect 2690 493 2697 496
rect 2694 426 2697 493
rect 2694 423 2701 426
rect 2590 313 2597 316
rect 2594 293 2597 313
rect 2546 283 2565 286
rect 2466 183 2469 206
rect 2370 123 2373 146
rect 2434 133 2437 176
rect 2450 133 2461 136
rect 2458 113 2461 126
rect 2466 103 2469 126
rect 2474 113 2477 126
rect 2482 113 2485 213
rect 2490 163 2493 206
rect 2522 193 2525 206
rect 2546 203 2549 216
rect 2490 133 2493 146
rect 2490 103 2493 116
rect 2506 103 2509 126
rect 2514 123 2517 136
rect 2530 133 2533 156
rect 2562 153 2565 283
rect 2586 193 2589 216
rect 2634 213 2637 326
rect 2642 213 2645 336
rect 2666 333 2677 336
rect 2682 316 2685 326
rect 2690 323 2693 416
rect 2698 316 2701 423
rect 2706 353 2709 513
rect 2714 333 2717 416
rect 2722 413 2725 516
rect 2730 403 2733 606
rect 2770 593 2773 616
rect 2818 566 2821 733
rect 2826 713 2829 726
rect 2810 563 2821 566
rect 2738 513 2741 536
rect 2778 533 2781 546
rect 2754 416 2757 526
rect 2786 513 2789 536
rect 2810 446 2813 563
rect 2810 443 2821 446
rect 2738 396 2741 416
rect 2746 403 2749 416
rect 2754 413 2765 416
rect 2754 396 2757 406
rect 2762 403 2765 413
rect 2650 303 2653 316
rect 2682 313 2701 316
rect 2714 313 2717 326
rect 2682 286 2685 313
rect 2682 283 2693 286
rect 2650 223 2653 246
rect 2674 203 2685 206
rect 2554 123 2557 146
rect 2674 133 2677 146
rect 2618 123 2629 126
rect 2626 113 2637 116
rect 2690 103 2693 283
rect 2722 276 2725 366
rect 2730 316 2733 396
rect 2738 393 2757 396
rect 2738 333 2741 386
rect 2730 313 2737 316
rect 2714 273 2725 276
rect 2698 213 2701 226
rect 2706 193 2709 206
rect 2714 203 2717 273
rect 2734 266 2737 313
rect 2746 303 2749 326
rect 2754 266 2757 356
rect 2730 263 2737 266
rect 2746 263 2757 266
rect 2730 203 2733 263
rect 2706 133 2709 156
rect 2722 133 2725 166
rect 2738 153 2741 216
rect 2746 203 2749 263
rect 2762 163 2765 226
rect 2786 223 2789 426
rect 2818 423 2821 443
rect 2834 436 2837 746
rect 2850 733 2853 923
rect 2866 826 2869 1076
rect 2874 1013 2877 1126
rect 2874 963 2877 1006
rect 2882 1003 2885 1146
rect 2890 1133 2893 1216
rect 2890 1113 2893 1126
rect 2890 996 2893 1026
rect 2882 993 2893 996
rect 2874 903 2877 926
rect 2882 913 2885 993
rect 2898 943 2901 1403
rect 2930 1396 2933 1443
rect 2922 1393 2933 1396
rect 2906 1223 2909 1316
rect 2906 1193 2909 1206
rect 2914 1203 2917 1336
rect 2922 1293 2925 1393
rect 2938 1343 2941 1536
rect 2954 1426 2957 1516
rect 2946 1423 2957 1426
rect 2946 1326 2949 1423
rect 2930 1313 2933 1326
rect 2938 1323 2949 1326
rect 2938 1306 2941 1323
rect 2930 1303 2941 1306
rect 2922 1186 2925 1216
rect 2930 1203 2933 1303
rect 2906 1183 2925 1186
rect 2906 1123 2909 1183
rect 2914 1133 2917 1176
rect 2922 1133 2925 1146
rect 2922 1103 2925 1126
rect 2906 993 2909 1016
rect 2914 983 2917 1006
rect 2922 973 2925 1096
rect 2938 1003 2941 1216
rect 2946 1193 2949 1206
rect 2946 1123 2949 1136
rect 2946 996 2949 1026
rect 2938 993 2949 996
rect 2890 923 2901 926
rect 2890 863 2893 906
rect 2898 903 2901 916
rect 2914 876 2917 936
rect 2906 873 2917 876
rect 2858 823 2869 826
rect 2858 793 2861 816
rect 2866 813 2869 823
rect 2866 783 2869 806
rect 2874 746 2877 816
rect 2890 813 2893 826
rect 2898 813 2901 836
rect 2906 813 2909 873
rect 2914 833 2917 866
rect 2898 793 2901 806
rect 2914 793 2917 826
rect 2922 823 2925 926
rect 2930 916 2933 946
rect 2938 933 2941 993
rect 2930 913 2937 916
rect 2934 846 2937 913
rect 2930 843 2937 846
rect 2922 803 2925 816
rect 2858 743 2877 746
rect 2850 703 2853 726
rect 2858 716 2861 743
rect 2866 733 2885 736
rect 2858 713 2865 716
rect 2842 603 2845 656
rect 2850 536 2853 696
rect 2862 646 2865 713
rect 2858 643 2865 646
rect 2858 613 2861 643
rect 2866 613 2869 626
rect 2858 543 2861 606
rect 2874 603 2877 726
rect 2882 613 2885 733
rect 2890 633 2893 716
rect 2898 713 2901 726
rect 2906 603 2909 736
rect 2914 733 2917 776
rect 2842 533 2853 536
rect 2874 533 2877 556
rect 2882 516 2885 536
rect 2914 533 2917 616
rect 2922 603 2925 786
rect 2930 733 2933 843
rect 2946 833 2949 986
rect 2954 953 2957 1416
rect 2962 1366 2965 1476
rect 2970 1383 2973 1553
rect 2986 1436 2989 1563
rect 2982 1433 2989 1436
rect 2982 1376 2985 1433
rect 3010 1426 3013 1626
rect 3010 1423 3021 1426
rect 2978 1373 2985 1376
rect 2962 1363 2969 1366
rect 2966 1286 2969 1363
rect 2978 1306 2981 1373
rect 2994 1343 2997 1406
rect 3002 1323 3005 1416
rect 3018 1316 3021 1423
rect 3010 1313 3021 1316
rect 2978 1303 2989 1306
rect 2966 1283 2973 1286
rect 2970 1176 2973 1283
rect 2966 1173 2973 1176
rect 2966 1026 2969 1173
rect 2986 1156 2989 1303
rect 2978 1153 2989 1156
rect 2978 1073 2981 1153
rect 3010 1136 3013 1313
rect 2994 1116 2997 1136
rect 3010 1133 3021 1136
rect 2990 1113 2997 1116
rect 2990 1036 2993 1113
rect 2990 1033 2997 1036
rect 2962 1023 2969 1026
rect 2962 943 2965 1023
rect 2994 1013 2997 1033
rect 2962 913 2965 926
rect 2970 903 2973 1006
rect 2986 926 2989 946
rect 2982 923 2989 926
rect 2938 813 2941 826
rect 2938 803 2949 806
rect 2954 803 2957 826
rect 2938 646 2941 726
rect 2962 656 2965 866
rect 2982 856 2985 923
rect 2994 863 2997 946
rect 3002 933 3005 1126
rect 3018 966 3021 1133
rect 3010 963 3021 966
rect 3010 943 3013 963
rect 2982 853 2989 856
rect 2970 773 2973 806
rect 2978 713 2981 816
rect 2986 783 2989 853
rect 2994 723 2997 746
rect 3002 723 3005 736
rect 2962 653 2973 656
rect 2938 643 2949 646
rect 2930 613 2933 626
rect 2938 613 2941 636
rect 2946 626 2949 643
rect 2946 623 2957 626
rect 2874 513 2885 516
rect 2874 446 2877 513
rect 2874 443 2885 446
rect 2826 433 2837 436
rect 2818 403 2821 416
rect 2810 323 2813 336
rect 2786 203 2789 216
rect 2826 193 2829 433
rect 2834 423 2861 426
rect 2834 413 2837 423
rect 2842 403 2845 416
rect 2866 323 2869 416
rect 2882 413 2885 443
rect 2882 383 2885 406
rect 2890 333 2893 526
rect 2906 503 2909 516
rect 2922 423 2925 596
rect 2938 553 2941 606
rect 2954 566 2957 623
rect 2946 563 2957 566
rect 2930 523 2933 546
rect 2946 543 2949 563
rect 2970 546 2973 653
rect 2970 543 2981 546
rect 2938 533 2957 536
rect 2938 503 2941 526
rect 2946 486 2949 526
rect 2942 483 2949 486
rect 2898 386 2901 406
rect 2906 403 2925 406
rect 2930 403 2933 416
rect 2942 406 2945 483
rect 2938 403 2945 406
rect 2954 403 2957 533
rect 2978 456 2981 543
rect 2962 453 2981 456
rect 2962 436 2965 453
rect 2962 433 2973 436
rect 2898 383 2909 386
rect 2874 313 2877 326
rect 2898 306 2901 366
rect 2906 313 2909 383
rect 2914 336 2917 396
rect 2922 373 2925 403
rect 2914 333 2925 336
rect 2914 313 2917 326
rect 2922 306 2925 333
rect 2930 313 2933 396
rect 2938 333 2941 403
rect 2962 393 2965 426
rect 2954 323 2957 386
rect 2970 363 2973 433
rect 2858 193 2861 216
rect 2746 123 2749 146
rect 2826 136 2829 146
rect 2810 133 2829 136
rect 2810 123 2813 133
rect 2834 123 2837 156
rect 2866 123 2869 306
rect 2898 303 2909 306
rect 2922 303 2933 306
rect 2890 203 2893 226
rect 2890 136 2893 196
rect 2882 133 2893 136
rect 2898 136 2901 206
rect 2906 183 2909 303
rect 2922 213 2925 226
rect 2898 133 2909 136
rect 2922 133 2925 146
rect 2882 103 2885 133
rect 2890 123 2901 126
rect 2906 116 2909 133
rect 2930 126 2933 303
rect 2938 296 2941 316
rect 2938 293 2949 296
rect 2946 226 2949 293
rect 2938 223 2949 226
rect 2938 203 2941 223
rect 2938 133 2941 146
rect 2970 133 2973 336
rect 2914 123 2925 126
rect 2930 123 2941 126
rect 2914 116 2917 123
rect 2898 113 2917 116
rect 2922 103 2925 116
rect 2970 103 2973 116
rect 3033 37 3053 3003
rect 3057 13 3077 3027
rect 3094 2862 3786 2867
rect 3113 2817 3753 2818
rect 3094 2813 3753 2817
rect 3094 2812 3118 2813
rect 3094 2732 3725 2737
rect 3094 2615 3120 2617
rect 3094 2612 3689 2615
rect 3115 2610 3689 2612
rect 3112 2537 3652 2539
rect 3094 2534 3652 2537
rect 3094 2532 3117 2534
rect 3094 2416 3104 2417
rect 3094 2412 3621 2416
rect 3099 2411 3621 2412
rect 3094 2362 3587 2367
rect 3094 2262 3553 2267
rect 3112 2187 3524 2188
rect 3094 2183 3524 2187
rect 3094 2182 3117 2183
rect 3106 2167 3495 2168
rect 3094 2163 3495 2167
rect 3094 2162 3111 2163
rect 3094 2142 3469 2147
rect 3115 2017 3442 2018
rect 3094 2013 3442 2017
rect 3094 2012 3120 2013
rect 3094 1932 3414 1937
rect 1697 -11 1702 0
rect -322 -681 -38 -676
rect -22 -16 1702 -11
rect -558 -743 -552 -737
rect -322 -743 -317 -681
rect -258 -743 -251 -736
rect -22 -743 -17 -16
rect 3094 -431 3099 1917
rect 2678 -436 3099 -431
rect 332 -719 578 -701
rect 2136 -707 2450 -692
rect 42 -743 48 -719
rect 642 -743 648 -719
rect 942 -743 948 -719
rect 1242 -743 1248 -719
rect 1542 -743 1548 -719
rect 1842 -743 1848 -719
rect 2441 -743 2450 -707
rect 2678 -743 2683 -436
rect 3409 -475 3414 1932
rect 2764 -480 3414 -475
rect 2764 -721 2769 -480
rect 3437 -527 3442 2013
rect 3065 -532 3442 -527
rect 2764 -726 2770 -721
rect 2742 -743 2748 -737
rect 2765 -743 2770 -726
rect 3042 -743 3048 -737
rect 3065 -743 3070 -532
rect 3464 -556 3469 2142
rect 3490 -515 3495 2163
rect 3519 -498 3524 2183
rect 3548 -413 3553 2262
rect 3582 -111 3587 2362
rect 3616 189 3621 2411
rect 3647 789 3652 2534
rect 3684 1089 3689 2610
rect 3720 1389 3725 2732
rect 3748 1689 3753 2813
rect 3781 1989 3786 2862
rect 3817 2589 3822 3059
rect 3849 2889 3854 3087
rect 3849 2884 3900 2889
rect 3894 2861 3900 2867
rect 3817 2584 3900 2589
rect 3894 2561 3900 2567
rect 3871 2244 3889 2561
rect 3781 1984 3900 1989
rect 3894 1961 3900 1967
rect 3748 1684 3900 1689
rect 3894 1661 3900 1667
rect 3720 1384 3900 1389
rect 3894 1361 3900 1367
rect 3684 1084 3900 1089
rect 3894 1061 3900 1067
rect 3647 784 3900 789
rect 3894 761 3900 767
rect 3871 448 3889 727
rect 3616 184 3900 189
rect 3894 161 3900 167
rect 3582 -116 3900 -111
rect 3894 -139 3900 -133
rect 3880 -413 3900 -411
rect 3548 -416 3900 -413
rect 3548 -418 3885 -416
rect 3894 -439 3900 -433
rect 3519 -503 3821 -498
rect 3490 -520 3670 -515
rect 3365 -561 3469 -556
rect 3342 -743 3348 -737
rect 3365 -743 3370 -561
rect 3642 -743 3648 -737
rect 3665 -743 3670 -520
rect 3816 -711 3821 -503
rect 3816 -716 3900 -711
rect 3894 -739 3900 -733
<< gv1 >>
rect -856 4015 -854 4017
rect -556 4015 -554 4017
rect -256 4015 -254 4017
rect 44 4015 46 4017
rect 1544 4015 1546 4017
rect 1844 4015 1846 4017
rect 2144 4015 2146 4017
rect 2444 4015 2446 4017
rect 2744 4015 2746 4017
rect 3344 4015 3346 4017
rect 3644 4015 3646 4017
rect 344 3982 346 3984
rect 644 3982 646 3984
rect 1244 3982 1246 3984
rect 945 3975 947 3977
rect 950 3975 952 3977
rect 955 3975 957 3977
rect 1181 3975 1183 3977
rect 1186 3975 1188 3977
rect 1191 3975 1193 3977
rect 3043 3975 3045 3977
rect 3048 3975 3050 3977
rect 3053 3975 3055 3977
rect 3274 3975 3276 3977
rect 3279 3975 3281 3977
rect 3284 3975 3286 3977
rect 945 3970 947 3972
rect 950 3970 952 3972
rect 955 3970 957 3972
rect 1181 3970 1183 3972
rect 1186 3970 1188 3972
rect 1191 3970 1193 3972
rect 3043 3970 3045 3972
rect 3048 3970 3050 3972
rect 3053 3970 3055 3972
rect 3274 3970 3276 3972
rect 3279 3970 3281 3972
rect 3284 3970 3286 3972
rect 945 3965 947 3967
rect 950 3965 952 3967
rect 955 3965 957 3967
rect 1181 3965 1183 3967
rect 1186 3965 1188 3967
rect 1191 3965 1193 3967
rect 3043 3965 3045 3967
rect 3048 3965 3050 3967
rect 3053 3965 3055 3967
rect 3274 3965 3276 3967
rect 3279 3965 3281 3967
rect 3284 3965 3286 3967
rect -860 3763 -858 3765
rect 3896 3763 3898 3765
rect -827 3463 -825 3465
rect 3896 3463 3898 3465
rect -827 3163 -825 3165
rect 3896 3163 3898 3165
rect 39 2942 41 2944
rect 44 2942 46 2944
rect 49 2942 51 2944
rect 54 2942 56 2944
rect 39 2937 41 2939
rect 44 2937 46 2939
rect 49 2937 51 2939
rect 54 2937 56 2939
rect 3034 2936 3036 2938
rect 3039 2936 3041 2938
rect 3044 2936 3046 2938
rect 3049 2936 3051 2938
rect 39 2932 41 2934
rect 44 2932 46 2934
rect 49 2932 51 2934
rect 54 2932 56 2934
rect 3034 2931 3036 2933
rect 3039 2931 3041 2933
rect 3044 2931 3046 2933
rect 3049 2931 3051 2933
rect 39 2927 41 2929
rect 44 2927 46 2929
rect 49 2927 51 2929
rect 54 2927 56 2929
rect 3034 2926 3036 2928
rect 3039 2926 3041 2928
rect 3044 2926 3046 2928
rect 3049 2926 3051 2928
rect 39 2922 41 2924
rect 44 2922 46 2924
rect 49 2922 51 2924
rect 54 2922 56 2924
rect 3034 2921 3036 2923
rect 3039 2921 3041 2923
rect 3044 2921 3046 2923
rect 3049 2921 3051 2923
rect 39 2917 41 2919
rect 44 2917 46 2919
rect 49 2917 51 2919
rect 54 2917 56 2919
rect 3034 2916 3036 2918
rect 3039 2916 3041 2918
rect 3044 2916 3046 2918
rect 3049 2916 3051 2918
rect 39 2912 41 2914
rect 44 2912 46 2914
rect 49 2912 51 2914
rect 54 2912 56 2914
rect 3034 2911 3036 2913
rect 3039 2911 3041 2913
rect 3044 2911 3046 2913
rect 3049 2911 3051 2913
rect 39 2907 41 2909
rect 44 2907 46 2909
rect 49 2907 51 2909
rect 54 2907 56 2909
rect 3034 2906 3036 2908
rect 3039 2906 3041 2908
rect 3044 2906 3046 2908
rect 3049 2906 3051 2908
rect 39 2902 41 2904
rect 44 2902 46 2904
rect 49 2902 51 2904
rect 54 2902 56 2904
rect 3034 2901 3036 2903
rect 3039 2901 3041 2903
rect 3044 2901 3046 2903
rect 3049 2901 3051 2903
rect 3034 2896 3036 2898
rect 3039 2896 3041 2898
rect 3044 2896 3046 2898
rect 3049 2896 3051 2898
rect -827 2863 -825 2865
rect 3896 2863 3898 2865
rect -849 2818 -847 2820
rect -844 2818 -842 2820
rect 3896 2563 3898 2565
rect 3874 2558 3876 2560
rect 3879 2558 3881 2560
rect 3884 2558 3886 2560
rect -849 2554 -847 2556
rect -844 2554 -842 2556
rect 3874 2553 3876 2555
rect 3879 2553 3881 2555
rect 3884 2553 3886 2555
rect -860 2511 -858 2513
rect 3874 2250 3876 2252
rect 3879 2250 3881 2252
rect 3884 2250 3886 2252
rect 3874 2245 3876 2247
rect 3879 2245 3881 2247
rect 3884 2245 3886 2247
rect -860 1963 -858 1965
rect 3896 1963 3898 1965
rect -860 1663 -858 1665
rect 3896 1663 3898 1665
rect -827 1363 -825 1365
rect 3896 1363 3898 1365
rect -827 1063 -825 1065
rect 3896 1063 3898 1065
rect -849 1027 -847 1029
rect -844 1027 -842 1029
rect 3896 763 3898 765
rect -849 757 -847 759
rect -844 757 -842 759
rect 3874 724 3876 726
rect 3879 724 3881 726
rect 3884 724 3886 726
rect 3874 719 3876 721
rect 3879 719 3881 721
rect 3884 719 3886 721
rect 3874 454 3876 456
rect 3879 454 3881 456
rect 3884 454 3886 456
rect 3874 449 3876 451
rect 3879 449 3881 451
rect 3884 449 3886 451
rect 39 432 41 434
rect 44 432 46 434
rect 49 432 51 434
rect 54 432 56 434
rect 39 427 41 429
rect 44 427 46 429
rect 49 427 51 429
rect 54 427 56 429
rect 39 422 41 424
rect 44 422 46 424
rect 49 422 51 424
rect 54 422 56 424
rect 39 417 41 419
rect 44 417 46 419
rect 49 417 51 419
rect 54 417 56 419
rect 39 412 41 414
rect 44 412 46 414
rect 49 412 51 414
rect 54 412 56 414
rect 39 407 41 409
rect 44 407 46 409
rect 49 407 51 409
rect 54 407 56 409
rect 39 402 41 404
rect 44 402 46 404
rect 49 402 51 404
rect 54 402 56 404
rect 39 397 41 399
rect 44 397 46 399
rect 49 397 51 399
rect 54 397 56 399
rect 39 392 41 394
rect 44 392 46 394
rect 49 392 51 394
rect 54 392 56 394
rect 3034 221 3036 223
rect 3039 221 3041 223
rect 3044 221 3046 223
rect 3049 221 3051 223
rect 3034 216 3036 218
rect 3039 216 3041 218
rect 3044 216 3046 218
rect 3049 216 3051 218
rect 3034 211 3036 213
rect 3039 211 3041 213
rect 3044 211 3046 213
rect 3049 211 3051 213
rect 3034 206 3036 208
rect 3039 206 3041 208
rect 3044 206 3046 208
rect 3049 206 3051 208
rect 3034 201 3036 203
rect 3039 201 3041 203
rect 3044 201 3046 203
rect 3049 201 3051 203
rect 3034 196 3036 198
rect 3039 196 3041 198
rect 3044 196 3046 198
rect 3049 196 3051 198
rect 3034 191 3036 193
rect 3039 191 3041 193
rect 3044 191 3046 193
rect 3049 191 3051 193
rect 3034 186 3036 188
rect 3039 186 3041 188
rect 3044 186 3046 188
rect 3049 186 3051 188
rect 3034 181 3036 183
rect 3039 181 3041 183
rect 3044 181 3046 183
rect 3049 181 3051 183
rect -860 163 -858 165
rect 3896 163 3898 165
rect -820 10 -818 12
rect -815 10 -813 12
rect -810 10 -808 12
rect -820 5 -818 7
rect -815 5 -813 7
rect -810 5 -808 7
rect -820 0 -818 2
rect -815 0 -813 2
rect -810 0 -808 2
rect -820 -75 -818 -73
rect -815 -75 -813 -73
rect -810 -75 -808 -73
rect -820 -80 -818 -78
rect -815 -80 -813 -78
rect -810 -80 -808 -78
rect -820 -85 -818 -83
rect -815 -85 -813 -83
rect -810 -85 -808 -83
rect -860 -137 -858 -135
rect 3896 -137 3898 -135
rect -860 -437 -858 -435
rect 3896 -437 3898 -435
rect 2137 -696 2139 -694
rect 2142 -696 2144 -694
rect 2442 -696 2444 -694
rect 2447 -696 2449 -694
rect 2137 -701 2139 -699
rect 2142 -701 2144 -699
rect 2442 -701 2444 -699
rect 2447 -701 2449 -699
rect 335 -706 337 -704
rect 340 -706 342 -704
rect 345 -706 347 -704
rect 563 -706 565 -704
rect 568 -706 570 -704
rect 573 -706 575 -704
rect 2137 -706 2139 -704
rect 2142 -706 2144 -704
rect 2442 -706 2444 -704
rect 2447 -706 2449 -704
rect 335 -711 337 -709
rect 340 -711 342 -709
rect 345 -711 347 -709
rect 563 -711 565 -709
rect 568 -711 570 -709
rect 573 -711 575 -709
rect 335 -716 337 -714
rect 340 -716 342 -714
rect 345 -716 347 -714
rect 563 -716 565 -714
rect 568 -716 570 -714
rect 573 -716 575 -714
rect 44 -723 46 -721
rect 644 -723 646 -721
rect 944 -723 946 -721
rect 1244 -723 1246 -721
rect 1544 -723 1546 -721
rect 1844 -723 1846 -721
rect -863 -731 -861 -729
rect 3896 -737 3898 -735
rect -850 -741 -848 -739
rect -556 -741 -554 -739
rect -256 -741 -254 -739
rect 2744 -741 2746 -739
rect 3044 -741 3046 -739
rect 3344 -741 3346 -739
rect 3644 -741 3646 -739
<< metal3 >>
rect 1849 3022 1886 3027
rect 2225 2992 2286 2997
rect 625 2982 710 2987
rect 625 2977 630 2982
rect 601 2972 630 2977
rect 705 2977 710 2982
rect 705 2972 750 2977
rect 1913 2972 2070 2977
rect 401 2962 502 2967
rect 521 2962 694 2967
rect 401 2957 406 2962
rect 321 2952 406 2957
rect 497 2957 502 2962
rect 497 2952 646 2957
rect 1801 2952 1910 2957
rect 529 2942 614 2947
rect 633 2942 670 2947
rect 945 2942 1014 2947
rect 1065 2942 1174 2947
rect 1297 2942 1318 2947
rect 1473 2942 1542 2947
rect 1681 2942 1726 2947
rect 417 2932 478 2937
rect 577 2932 766 2937
rect 81 2922 126 2927
rect 313 2922 518 2927
rect 545 2922 574 2927
rect 649 2922 702 2927
rect 745 2922 798 2927
rect 1145 2922 1462 2927
rect 545 2917 550 2922
rect 1457 2917 1462 2922
rect 1553 2922 1654 2927
rect 1673 2922 1710 2927
rect 1921 2922 1926 2967
rect 2761 2952 2838 2957
rect 2761 2947 2766 2952
rect 2049 2942 2094 2947
rect 2209 2942 2270 2947
rect 2313 2942 2766 2947
rect 2833 2947 2838 2952
rect 2897 2952 2934 2957
rect 2897 2947 2902 2952
rect 2833 2942 2902 2947
rect 2913 2942 2958 2947
rect 2033 2932 2198 2937
rect 2777 2932 2822 2937
rect 2857 2922 2886 2927
rect 1553 2917 1558 2922
rect 241 2912 550 2917
rect 561 2912 598 2917
rect 737 2912 790 2917
rect 889 2912 990 2917
rect 1113 2912 1166 2917
rect 1457 2912 1558 2917
rect 1649 2917 1654 2922
rect 1649 2912 1774 2917
rect 2177 2912 2206 2917
rect 265 2902 358 2907
rect 505 2902 566 2907
rect 2049 2902 2166 2907
rect 337 2882 390 2887
rect 729 2882 758 2887
rect 1689 2882 1718 2887
rect 3093 2867 3100 2868
rect 1457 2862 1502 2867
rect 2905 2862 3100 2867
rect 3093 2861 3100 2862
rect 425 2852 646 2857
rect 2065 2852 2174 2857
rect 2689 2852 2766 2857
rect 169 2842 214 2847
rect 425 2837 430 2852
rect 177 2832 294 2837
rect 401 2832 430 2837
rect 641 2837 646 2852
rect 777 2842 822 2847
rect 1089 2842 1150 2847
rect 1209 2842 1342 2847
rect 1561 2842 1670 2847
rect 1561 2837 1566 2842
rect 641 2832 670 2837
rect 761 2832 822 2837
rect 1009 2832 1062 2837
rect 1105 2832 1222 2837
rect 1361 2832 1414 2837
rect 1505 2832 1566 2837
rect 1665 2837 1670 2842
rect 2257 2842 2366 2847
rect 2257 2837 2262 2842
rect 1665 2832 2086 2837
rect 2081 2827 2086 2832
rect 2145 2832 2262 2837
rect 2361 2837 2366 2842
rect 2473 2842 2590 2847
rect 2473 2837 2478 2842
rect 2361 2832 2478 2837
rect 2585 2837 2590 2842
rect 2633 2837 2750 2842
rect 2585 2832 2638 2837
rect 2745 2832 2830 2837
rect 2145 2827 2150 2832
rect 129 2822 166 2827
rect 369 2822 398 2827
rect 409 2822 454 2827
rect 505 2822 558 2827
rect 633 2822 750 2827
rect 785 2822 838 2827
rect 897 2822 998 2827
rect 1201 2822 1238 2827
rect 1617 2822 1638 2827
rect 2081 2822 2150 2827
rect 2169 2822 2342 2827
rect 145 2812 206 2817
rect 497 2812 526 2817
rect 537 2812 582 2817
rect 593 2812 622 2817
rect 793 2812 846 2817
rect 1001 2812 1030 2817
rect 1057 2812 1086 2817
rect 1193 2812 1246 2817
rect 1561 2812 1654 2817
rect 2193 2812 2222 2817
rect 2329 2812 2462 2817
rect 2521 2812 2550 2817
rect 2217 2807 2334 2812
rect 121 2802 302 2807
rect 313 2802 342 2807
rect 457 2802 622 2807
rect 1065 2802 1142 2807
rect 1305 2802 1374 2807
rect 1465 2802 1494 2807
rect 1609 2802 1670 2807
rect 1697 2802 1766 2807
rect 2409 2802 2478 2807
rect 2577 2802 2582 2827
rect 2657 2822 2870 2827
rect 2889 2822 3014 2827
rect 3009 2817 3014 2822
rect 3093 2817 3100 2818
rect 2593 2812 2638 2817
rect 2689 2812 2710 2817
rect 2825 2812 2902 2817
rect 3009 2812 3100 2817
rect 3093 2811 3100 2812
rect 2705 2802 2734 2807
rect 2705 2797 2710 2802
rect 233 2792 262 2797
rect 257 2787 262 2792
rect 337 2792 366 2797
rect 529 2792 638 2797
rect 953 2792 1062 2797
rect 1153 2792 1182 2797
rect 1289 2792 1326 2797
rect 1577 2792 2030 2797
rect 2057 2792 2126 2797
rect 2233 2792 2294 2797
rect 2457 2792 2558 2797
rect 2633 2792 2710 2797
rect 2857 2792 2958 2797
rect 337 2787 342 2792
rect 257 2782 342 2787
rect 561 2782 742 2787
rect 1041 2782 1070 2787
rect 1065 2777 1070 2782
rect 1145 2782 1302 2787
rect 1329 2782 1374 2787
rect 1705 2782 1822 2787
rect 2625 2782 2654 2787
rect 1145 2777 1150 2782
rect 537 2772 574 2777
rect 825 2772 990 2777
rect 1065 2772 1150 2777
rect 1169 2772 1342 2777
rect 1641 2772 1718 2777
rect 2649 2772 2710 2777
rect 1233 2762 1254 2767
rect 1529 2762 1582 2767
rect 2433 2762 2462 2767
rect 2553 2762 2838 2767
rect 113 2752 190 2757
rect 241 2752 350 2757
rect 361 2752 390 2757
rect 401 2752 542 2757
rect 1185 2752 1270 2757
rect 1905 2752 1926 2757
rect 2033 2752 2078 2757
rect 2537 2752 2630 2757
rect 169 2732 246 2737
rect 273 2727 278 2747
rect 377 2742 422 2747
rect 721 2742 742 2747
rect 753 2742 814 2747
rect 881 2742 1046 2747
rect 1065 2742 1134 2747
rect 1041 2737 1046 2742
rect 1233 2737 1238 2747
rect 1801 2742 1838 2747
rect 1929 2742 2142 2747
rect 2281 2742 2326 2747
rect 2377 2742 2510 2747
rect 2633 2742 2718 2747
rect 2833 2742 2870 2747
rect 2897 2742 2958 2747
rect 3093 2737 3100 2738
rect 345 2732 374 2737
rect 385 2732 566 2737
rect 577 2732 686 2737
rect 945 2732 1022 2737
rect 1041 2732 1142 2737
rect 1233 2732 1294 2737
rect 1665 2732 1774 2737
rect 1881 2732 1918 2737
rect 1969 2732 2030 2737
rect 2481 2732 2542 2737
rect 2617 2732 2678 2737
rect 3009 2732 3100 2737
rect 2257 2727 2358 2732
rect 3093 2731 3100 2732
rect 185 2722 310 2727
rect 329 2722 358 2727
rect 449 2722 558 2727
rect 705 2722 798 2727
rect 809 2722 854 2727
rect 1145 2722 1166 2727
rect 1369 2722 1438 2727
rect 1489 2722 1526 2727
rect 1761 2722 1870 2727
rect 2017 2722 2046 2727
rect 2233 2722 2262 2727
rect 2353 2722 2382 2727
rect 2465 2722 2542 2727
rect 2857 2722 2886 2727
rect 353 2717 454 2722
rect 1369 2717 1374 2722
rect 153 2712 182 2717
rect 561 2712 1014 2717
rect 1009 2707 1014 2712
rect 1177 2712 1374 2717
rect 1433 2717 1438 2722
rect 1865 2717 2006 2722
rect 1433 2712 1542 2717
rect 1657 2712 1718 2717
rect 1745 2712 1782 2717
rect 2001 2712 2278 2717
rect 2313 2712 2358 2717
rect 2489 2712 2854 2717
rect 2913 2712 3014 2717
rect 1177 2707 1182 2712
rect 81 2702 278 2707
rect 289 2702 342 2707
rect 361 2702 454 2707
rect 489 2702 558 2707
rect 657 2702 774 2707
rect 841 2702 870 2707
rect 1009 2702 1182 2707
rect 1873 2702 1982 2707
rect 2313 2702 2486 2707
rect 2505 2702 2654 2707
rect 1873 2697 1878 2702
rect 1977 2697 2126 2702
rect 209 2692 286 2697
rect 313 2692 494 2697
rect 721 2692 742 2697
rect 1385 2692 1422 2697
rect 1641 2692 1686 2697
rect 1697 2692 1878 2697
rect 2121 2692 2206 2697
rect 2369 2692 2478 2697
rect 2561 2692 2670 2697
rect 2473 2687 2566 2692
rect 2665 2687 2670 2692
rect 2809 2692 2838 2697
rect 2809 2687 2814 2692
rect 137 2682 166 2687
rect 385 2682 510 2687
rect 889 2682 990 2687
rect 161 2677 166 2682
rect 249 2677 390 2682
rect 889 2677 894 2682
rect 161 2672 254 2677
rect 409 2672 446 2677
rect 529 2672 702 2677
rect 529 2667 534 2672
rect 273 2662 398 2667
rect 457 2662 534 2667
rect 697 2667 702 2672
rect 833 2672 894 2677
rect 985 2677 990 2682
rect 1257 2682 1366 2687
rect 1889 2682 2110 2687
rect 2233 2682 2310 2687
rect 2585 2682 2646 2687
rect 2665 2682 2814 2687
rect 1257 2677 1262 2682
rect 985 2672 1262 2677
rect 1361 2677 1366 2682
rect 2105 2677 2238 2682
rect 1361 2672 1406 2677
rect 1713 2672 1742 2677
rect 1777 2672 2086 2677
rect 2473 2672 2566 2677
rect 833 2667 838 2672
rect 2281 2667 2390 2672
rect 2473 2667 2478 2672
rect 697 2662 838 2667
rect 857 2662 974 2667
rect 1281 2662 1342 2667
rect 2089 2662 2286 2667
rect 2385 2662 2478 2667
rect 2561 2667 2566 2672
rect 2561 2662 2606 2667
rect 393 2657 462 2662
rect 1737 2657 1966 2662
rect 601 2652 678 2657
rect 1273 2652 1390 2657
rect 1713 2652 1742 2657
rect 1961 2652 1990 2657
rect 2009 2652 2158 2657
rect 2297 2652 2374 2657
rect 2489 2652 2870 2657
rect 601 2647 606 2652
rect 353 2642 606 2647
rect 673 2647 678 2652
rect 1713 2647 1718 2652
rect 673 2642 758 2647
rect 1265 2642 1302 2647
rect 1553 2642 1718 2647
rect 1769 2642 1822 2647
rect 1841 2642 2238 2647
rect 2329 2642 2438 2647
rect 2553 2642 2614 2647
rect 617 2632 670 2637
rect 1153 2632 1222 2637
rect 1265 2632 1358 2637
rect 1801 2632 1950 2637
rect 1961 2632 2038 2637
rect 2057 2632 2078 2637
rect 2113 2632 2166 2637
rect 2281 2632 2342 2637
rect 2353 2632 2390 2637
rect 2417 2632 2710 2637
rect 2337 2627 2342 2632
rect 2417 2627 2422 2632
rect 177 2622 214 2627
rect 273 2622 302 2627
rect 401 2622 446 2627
rect 1145 2622 1190 2627
rect 1441 2622 1486 2627
rect 1729 2622 1822 2627
rect 1977 2622 2078 2627
rect 2097 2622 2126 2627
rect 313 2612 390 2617
rect 457 2612 534 2617
rect 721 2612 822 2617
rect 1017 2612 1094 2617
rect 1137 2612 1182 2617
rect 1449 2612 1494 2617
rect 1585 2612 1702 2617
rect 1713 2612 1894 2617
rect 2017 2612 2070 2617
rect 2145 2612 2262 2617
rect 385 2607 462 2612
rect 1713 2607 1718 2612
rect 2145 2607 2150 2612
rect 337 2602 358 2607
rect 1001 2602 1158 2607
rect 1241 2602 1350 2607
rect 1553 2602 1718 2607
rect 1729 2602 1782 2607
rect 1825 2602 1982 2607
rect 1993 2602 2150 2607
rect 1553 2597 1558 2602
rect 1729 2597 1734 2602
rect 2257 2597 2262 2612
rect 2321 2607 2326 2627
rect 2337 2622 2422 2627
rect 2433 2622 2462 2627
rect 2457 2617 2462 2622
rect 2569 2622 2678 2627
rect 2569 2617 2574 2622
rect 3093 2617 3100 2618
rect 2457 2612 2574 2617
rect 2681 2612 2798 2617
rect 2913 2612 3100 2617
rect 3093 2611 3100 2612
rect 2273 2602 2326 2607
rect 2345 2602 2382 2607
rect 2737 2602 2782 2607
rect 129 2592 206 2597
rect 217 2592 270 2597
rect 345 2592 422 2597
rect 577 2592 630 2597
rect 769 2592 838 2597
rect 929 2592 974 2597
rect 1065 2592 1206 2597
rect 1225 2592 1262 2597
rect 1377 2592 1558 2597
rect 1569 2592 1614 2597
rect 1681 2592 1734 2597
rect 1793 2592 1910 2597
rect 1921 2592 2126 2597
rect 2153 2592 2206 2597
rect 2257 2592 2422 2597
rect 2593 2592 2622 2597
rect 2673 2592 2830 2597
rect 2873 2592 2958 2597
rect 185 2582 302 2587
rect 409 2582 646 2587
rect 857 2582 1318 2587
rect 1361 2582 1438 2587
rect 1537 2582 1566 2587
rect 1625 2582 1726 2587
rect 1769 2582 1830 2587
rect 2033 2582 2182 2587
rect 2257 2582 2286 2587
rect 2305 2582 2406 2587
rect 1361 2577 1366 2582
rect 1561 2577 1630 2582
rect 2257 2577 2262 2582
rect 793 2572 846 2577
rect 841 2567 846 2572
rect 929 2572 958 2577
rect 1041 2572 1246 2577
rect 1337 2572 1366 2577
rect 1385 2572 1526 2577
rect 929 2567 934 2572
rect 1241 2567 1342 2572
rect 1521 2567 1526 2572
rect 1673 2572 2014 2577
rect 1673 2567 1678 2572
rect 2009 2567 2014 2572
rect 2113 2572 2262 2577
rect 2289 2572 2318 2577
rect 2681 2572 2726 2577
rect 2113 2567 2118 2572
rect 841 2562 934 2567
rect 1521 2562 1678 2567
rect 1697 2562 1838 2567
rect 1849 2562 1934 2567
rect 2009 2562 2118 2567
rect 2145 2562 2246 2567
rect 2257 2562 2366 2567
rect 1113 2557 1222 2562
rect 617 2552 662 2557
rect 1089 2552 1118 2557
rect 1217 2552 1358 2557
rect 1905 2552 1950 2557
rect 2241 2552 2766 2557
rect 129 2542 206 2547
rect 385 2542 614 2547
rect 841 2542 982 2547
rect 1153 2542 1206 2547
rect 1321 2542 1382 2547
rect 1409 2542 1550 2547
rect 1569 2542 1614 2547
rect 1745 2542 1790 2547
rect 1889 2542 1918 2547
rect 1937 2542 1990 2547
rect 2137 2542 2246 2547
rect 2433 2542 2630 2547
rect 2721 2542 2790 2547
rect 2897 2542 2958 2547
rect 1409 2537 1414 2542
rect 193 2532 246 2537
rect 521 2532 670 2537
rect 705 2532 734 2537
rect 1009 2532 1222 2537
rect 1265 2532 1294 2537
rect 1385 2532 1414 2537
rect 1545 2537 1550 2542
rect 2241 2537 2438 2542
rect 3093 2537 3100 2538
rect 1545 2532 1622 2537
rect 1841 2532 1958 2537
rect 1977 2532 2110 2537
rect 2457 2532 2494 2537
rect 2585 2532 2694 2537
rect 3009 2532 3100 2537
rect 753 2527 854 2532
rect 1289 2527 1390 2532
rect 3093 2531 3100 2532
rect 81 2522 158 2527
rect 609 2522 654 2527
rect 665 2522 758 2527
rect 849 2522 1054 2527
rect 1097 2522 1214 2527
rect 217 2517 294 2522
rect 1425 2517 1430 2527
rect 1481 2522 1526 2527
rect 1537 2522 1662 2527
rect 1721 2522 1870 2527
rect 1889 2522 2046 2527
rect 2241 2522 2358 2527
rect 2513 2522 2550 2527
rect 2713 2522 2838 2527
rect 2913 2522 3006 2527
rect 193 2512 222 2517
rect 289 2512 406 2517
rect 713 2512 846 2517
rect 865 2512 894 2517
rect 865 2507 870 2512
rect 113 2502 214 2507
rect 249 2502 278 2507
rect 273 2487 278 2502
rect 417 2502 526 2507
rect 833 2502 870 2507
rect 417 2487 422 2502
rect 889 2497 894 2512
rect 1049 2512 1182 2517
rect 1313 2512 1334 2517
rect 1425 2512 1518 2517
rect 1681 2512 1726 2517
rect 1049 2497 1054 2512
rect 1425 2507 1430 2512
rect 1073 2502 1430 2507
rect 1553 2502 1854 2507
rect 1953 2502 2142 2507
rect 2153 2502 2214 2507
rect 2313 2502 2374 2507
rect 2745 2502 2854 2507
rect 889 2492 1054 2497
rect 1665 2492 2022 2497
rect 2033 2492 2078 2497
rect 2097 2492 2406 2497
rect 2401 2487 2406 2492
rect 273 2482 422 2487
rect 1977 2482 2390 2487
rect 2401 2482 2478 2487
rect 1745 2477 1902 2482
rect 1169 2472 1534 2477
rect 1553 2472 1574 2477
rect 1593 2472 1702 2477
rect 1721 2472 1750 2477
rect 1897 2472 2118 2477
rect 2497 2472 2582 2477
rect 1169 2467 1174 2472
rect 593 2462 854 2467
rect 961 2462 1174 2467
rect 1529 2467 1534 2472
rect 1593 2467 1598 2472
rect 1529 2462 1598 2467
rect 1697 2467 1702 2472
rect 2225 2467 2502 2472
rect 2577 2467 2582 2472
rect 1697 2462 1886 2467
rect 2041 2462 2230 2467
rect 2577 2462 2670 2467
rect 593 2447 598 2462
rect 849 2457 854 2462
rect 849 2452 942 2457
rect 249 2442 278 2447
rect 569 2442 598 2447
rect 937 2447 942 2452
rect 1201 2452 1286 2457
rect 1353 2452 1758 2457
rect 1873 2452 2102 2457
rect 2121 2452 2150 2457
rect 2241 2452 2566 2457
rect 1201 2447 1206 2452
rect 937 2442 1054 2447
rect 1049 2437 1054 2442
rect 1185 2442 1206 2447
rect 1281 2447 1286 2452
rect 1873 2447 1878 2452
rect 2145 2447 2246 2452
rect 1281 2442 1310 2447
rect 1569 2442 1814 2447
rect 1825 2442 1878 2447
rect 1897 2442 1934 2447
rect 2265 2442 2422 2447
rect 2449 2442 2494 2447
rect 1185 2437 1190 2442
rect 1825 2437 1830 2442
rect 217 2432 326 2437
rect 377 2432 494 2437
rect 529 2432 718 2437
rect 729 2432 838 2437
rect 1049 2432 1190 2437
rect 1209 2432 1270 2437
rect 1545 2432 1830 2437
rect 1841 2432 1870 2437
rect 1905 2432 2318 2437
rect 2425 2432 2470 2437
rect 2617 2432 2694 2437
rect 1905 2427 1910 2432
rect 2617 2427 2622 2432
rect 313 2422 342 2427
rect 545 2422 590 2427
rect 737 2422 902 2427
rect 921 2422 1030 2427
rect 1329 2422 1542 2427
rect 1585 2422 1646 2427
rect 1713 2422 1742 2427
rect 1809 2422 1910 2427
rect 2361 2422 2622 2427
rect 2689 2427 2694 2432
rect 2689 2422 2742 2427
rect 2913 2422 3014 2427
rect 1929 2417 2190 2422
rect 257 2412 294 2417
rect 305 2412 358 2417
rect 705 2412 798 2417
rect 865 2412 902 2417
rect 1441 2412 1470 2417
rect 1465 2407 1470 2412
rect 1545 2412 1678 2417
rect 1705 2412 1750 2417
rect 1785 2412 1934 2417
rect 2185 2412 2214 2417
rect 2313 2412 2406 2417
rect 2641 2412 2678 2417
rect 1545 2407 1550 2412
rect 2209 2407 2214 2412
rect 2705 2407 2710 2422
rect 3009 2417 3014 2422
rect 3093 2417 3100 2418
rect 3009 2412 3100 2417
rect 3093 2411 3100 2412
rect 129 2402 190 2407
rect 273 2402 342 2407
rect 369 2402 454 2407
rect 769 2402 870 2407
rect 985 2402 1030 2407
rect 1465 2402 1550 2407
rect 1889 2402 2190 2407
rect 2209 2402 2318 2407
rect 2313 2397 2318 2402
rect 2433 2402 2486 2407
rect 2633 2402 2654 2407
rect 2705 2402 2734 2407
rect 2433 2397 2438 2402
rect 193 2392 214 2397
rect 241 2392 262 2397
rect 281 2392 390 2397
rect 681 2392 766 2397
rect 953 2392 982 2397
rect 1145 2392 1214 2397
rect 1345 2392 1446 2397
rect 1601 2392 1670 2397
rect 1873 2392 1942 2397
rect 2073 2392 2118 2397
rect 2129 2392 2166 2397
rect 2313 2392 2438 2397
rect 2457 2392 2558 2397
rect 2569 2392 2782 2397
rect 2801 2392 2894 2397
rect 2913 2392 2958 2397
rect 1977 2387 2054 2392
rect 2129 2387 2134 2392
rect 329 2382 470 2387
rect 641 2382 710 2387
rect 889 2382 918 2387
rect 993 2382 1262 2387
rect 1297 2382 1566 2387
rect 1913 2382 1982 2387
rect 2049 2382 2134 2387
rect 2169 2382 2230 2387
rect 2593 2382 2726 2387
rect 913 2377 998 2382
rect 233 2372 318 2377
rect -6 2367 1 2368
rect 313 2367 318 2372
rect 377 2372 406 2377
rect 1177 2372 1246 2377
rect 1305 2372 1406 2377
rect 1993 2372 2294 2377
rect 2569 2372 2598 2377
rect 377 2367 382 2372
rect 1057 2367 1158 2372
rect 2593 2367 2598 2372
rect 2665 2372 2718 2377
rect 2665 2367 2670 2372
rect 3093 2367 3100 2368
rect -6 2362 70 2367
rect 257 2362 278 2367
rect 313 2362 382 2367
rect 1033 2362 1062 2367
rect 1153 2362 1430 2367
rect 1585 2362 1614 2367
rect 1969 2362 2006 2367
rect 2129 2362 2158 2367
rect 2257 2362 2286 2367
rect 2593 2362 2670 2367
rect 2689 2362 2750 2367
rect 2881 2362 3100 2367
rect -6 2361 1 2362
rect 2153 2357 2262 2362
rect 3093 2361 3100 2362
rect 65 2352 174 2357
rect 833 2352 918 2357
rect 1081 2352 1206 2357
rect 1233 2352 1318 2357
rect 2769 2352 2862 2357
rect 833 2347 838 2352
rect 241 2342 366 2347
rect 393 2342 502 2347
rect 697 2342 726 2347
rect 809 2342 838 2347
rect 913 2347 918 2352
rect 2769 2347 2774 2352
rect 913 2342 942 2347
rect 1017 2342 1070 2347
rect 1289 2342 1390 2347
rect 1745 2342 1806 2347
rect 1825 2342 1870 2347
rect 553 2332 614 2337
rect 817 2332 870 2337
rect 1089 2332 1206 2337
rect 1537 2332 1558 2337
rect 1585 2332 1662 2337
rect 305 2327 422 2332
rect 1089 2327 1094 2332
rect 201 2322 262 2327
rect 281 2322 310 2327
rect 417 2322 446 2327
rect 825 2322 1094 2327
rect 1201 2327 1206 2332
rect 1585 2327 1590 2332
rect 1201 2322 1246 2327
rect 1561 2322 1590 2327
rect 1657 2327 1662 2332
rect 1881 2327 1886 2347
rect 1977 2342 2214 2347
rect 2657 2342 2710 2347
rect 2737 2342 2774 2347
rect 2857 2347 2862 2352
rect 2857 2342 2902 2347
rect 2321 2332 2390 2337
rect 2321 2327 2326 2332
rect 1657 2322 1686 2327
rect 1881 2322 2118 2327
rect 2113 2317 2118 2322
rect 2225 2322 2326 2327
rect 2385 2327 2390 2332
rect 2617 2327 2686 2332
rect 2385 2322 2622 2327
rect 2681 2322 2934 2327
rect 2225 2317 2230 2322
rect 217 2312 326 2317
rect 353 2312 406 2317
rect 449 2312 478 2317
rect 569 2312 678 2317
rect 689 2312 806 2317
rect 129 2302 198 2307
rect 353 2302 358 2312
rect 689 2307 694 2312
rect 385 2302 422 2307
rect 665 2302 694 2307
rect 801 2307 806 2312
rect 921 2312 1222 2317
rect 1297 2312 1326 2317
rect 1593 2312 1622 2317
rect 1729 2312 1782 2317
rect 2113 2312 2230 2317
rect 2633 2312 2662 2317
rect 921 2307 926 2312
rect 801 2302 926 2307
rect 945 2302 1006 2307
rect 1105 2302 1126 2307
rect 1425 2302 1718 2307
rect 1793 2302 1822 2307
rect 1897 2302 1998 2307
rect 2041 2302 2094 2307
rect 2337 2302 2374 2307
rect 2457 2302 2478 2307
rect 2697 2302 2734 2307
rect 2873 2302 2918 2307
rect -6 2297 1 2298
rect 1105 2297 1110 2302
rect 1713 2297 1798 2302
rect -6 2292 70 2297
rect 401 2292 542 2297
rect 985 2292 1110 2297
rect 1249 2292 1318 2297
rect 2409 2292 2598 2297
rect -6 2291 1 2292
rect 1617 2287 1686 2292
rect 257 2282 334 2287
rect 561 2282 662 2287
rect 1105 2282 1622 2287
rect 1681 2282 2054 2287
rect 2073 2282 2102 2287
rect 257 2277 262 2282
rect 329 2277 566 2282
rect 657 2277 662 2282
rect 113 2272 262 2277
rect 657 2272 686 2277
rect 1633 2272 1670 2277
rect 2137 2272 2174 2277
rect 2193 2272 2390 2277
rect 2009 2267 2118 2272
rect 2193 2267 2198 2272
rect 329 2262 702 2267
rect 721 2262 1054 2267
rect 721 2257 726 2262
rect 273 2252 510 2257
rect 505 2247 510 2252
rect 681 2252 726 2257
rect 1049 2257 1054 2262
rect 1481 2262 1606 2267
rect 1481 2257 1486 2262
rect 1049 2252 1078 2257
rect 1161 2252 1350 2257
rect 1457 2252 1486 2257
rect 1601 2257 1606 2262
rect 1697 2262 2014 2267
rect 2113 2262 2198 2267
rect 2385 2267 2390 2272
rect 2409 2272 2478 2277
rect 2409 2267 2414 2272
rect 2385 2262 2414 2267
rect 2473 2267 2478 2272
rect 3093 2267 3100 2268
rect 2473 2262 2670 2267
rect 3009 2262 3100 2267
rect 1697 2257 1702 2262
rect 3093 2261 3100 2262
rect 1601 2252 1702 2257
rect 2025 2252 2126 2257
rect 2425 2252 2462 2257
rect 2729 2252 2822 2257
rect 681 2247 686 2252
rect 1913 2247 2030 2252
rect 2729 2247 2734 2252
rect 289 2242 422 2247
rect 465 2242 486 2247
rect 505 2242 686 2247
rect 705 2242 758 2247
rect 777 2242 798 2247
rect 1449 2242 1590 2247
rect 1585 2237 1590 2242
rect 1713 2242 1918 2247
rect 2049 2242 2414 2247
rect 1713 2237 1718 2242
rect 2409 2237 2414 2242
rect 2473 2242 2734 2247
rect 2817 2247 2822 2252
rect 2817 2242 2902 2247
rect 2473 2237 2478 2242
rect 377 2232 446 2237
rect 841 2232 1030 2237
rect 1057 2232 1166 2237
rect 1305 2232 1326 2237
rect 1481 2232 1510 2237
rect 1585 2232 1718 2237
rect 1937 2232 2054 2237
rect 2121 2232 2182 2237
rect 2409 2232 2478 2237
rect 2513 2232 2542 2237
rect 2609 2232 2742 2237
rect 345 2222 390 2227
rect 425 2222 630 2227
rect 681 2222 806 2227
rect 865 2222 910 2227
rect 1009 2222 1094 2227
rect 625 2212 630 2222
rect 1121 2217 1126 2227
rect 1265 2222 1302 2227
rect 1321 2222 1398 2227
rect 1473 2222 1550 2227
rect 2577 2222 2638 2227
rect 2665 2222 2806 2227
rect 697 2212 750 2217
rect 881 2212 926 2217
rect 937 2212 982 2217
rect 1001 2212 1126 2217
rect 1201 2212 1278 2217
rect 1337 2212 1382 2217
rect 1489 2212 1510 2217
rect 1745 2212 1766 2217
rect 1777 2212 1870 2217
rect 2001 2212 2326 2217
rect 2353 2212 2454 2217
rect 2561 2212 2606 2217
rect 2617 2212 2678 2217
rect 2689 2212 2710 2217
rect 2721 2212 2790 2217
rect 529 2202 742 2207
rect 793 2202 902 2207
rect 969 2202 998 2207
rect 737 2197 742 2202
rect 993 2197 998 2202
rect 1089 2202 1222 2207
rect 1641 2202 1726 2207
rect 1089 2197 1094 2202
rect 1641 2197 1646 2202
rect 153 2192 214 2197
rect 233 2192 294 2197
rect 321 2192 454 2197
rect 481 2192 566 2197
rect 609 2192 718 2197
rect 737 2192 950 2197
rect 993 2192 1094 2197
rect 1137 2192 1198 2197
rect 1225 2192 1278 2197
rect 1369 2192 1438 2197
rect 1481 2192 1518 2197
rect 1529 2192 1646 2197
rect 1721 2197 1726 2202
rect 2177 2202 2262 2207
rect 2649 2202 2718 2207
rect 2177 2197 2182 2202
rect 1721 2192 1750 2197
rect 1761 2192 1814 2197
rect 1913 2192 2182 2197
rect 2193 2192 2390 2197
rect 2449 2192 2566 2197
rect 2657 2192 2726 2197
rect 2833 2192 2838 2242
rect 2897 2237 2902 2242
rect 2897 2232 2974 2237
rect 2865 2192 2926 2197
rect 2993 2192 3070 2197
rect 209 2177 214 2192
rect 1745 2187 1750 2192
rect 2993 2187 2998 2192
rect 313 2182 342 2187
rect 785 2182 870 2187
rect 1113 2182 1174 2187
rect 1393 2182 1438 2187
rect 1641 2182 1726 2187
rect 1745 2182 1902 2187
rect 2145 2182 2214 2187
rect 2921 2182 2998 2187
rect 3065 2187 3070 2192
rect 3093 2187 3100 2188
rect 3065 2182 3100 2187
rect 313 2177 318 2182
rect 889 2177 998 2182
rect 1433 2177 1558 2182
rect 1641 2177 1646 2182
rect 1897 2177 1982 2182
rect 2145 2177 2150 2182
rect 3093 2181 3100 2182
rect 209 2172 318 2177
rect 449 2172 678 2177
rect 713 2172 894 2177
rect 993 2172 1414 2177
rect 1553 2172 1646 2177
rect 1825 2172 1862 2177
rect 1977 2172 2150 2177
rect 2289 2172 2462 2177
rect 2489 2172 2534 2177
rect 3093 2167 3100 2168
rect 465 2162 494 2167
rect 641 2162 710 2167
rect 745 2162 806 2167
rect 905 2162 982 2167
rect 1105 2162 1142 2167
rect 1513 2162 1534 2167
rect 1665 2162 1734 2167
rect 1857 2162 1958 2167
rect 2521 2162 2550 2167
rect 2857 2162 2918 2167
rect 3009 2162 3100 2167
rect 489 2157 494 2162
rect 561 2157 646 2162
rect 3093 2161 3100 2162
rect 489 2152 566 2157
rect 665 2152 958 2157
rect 1017 2152 1086 2157
rect 1273 2152 1358 2157
rect 1401 2152 1702 2157
rect 1713 2152 1798 2157
rect 1849 2152 1966 2157
rect 2033 2152 2374 2157
rect 2553 2152 2598 2157
rect 2705 2152 2734 2157
rect 2785 2152 2950 2157
rect 385 2142 430 2147
rect 585 2142 614 2147
rect 737 2142 798 2147
rect 841 2142 870 2147
rect 865 2137 870 2142
rect 961 2142 1046 2147
rect 1193 2142 1230 2147
rect 1329 2142 1374 2147
rect 1449 2142 1494 2147
rect 1793 2142 1830 2147
rect 1905 2142 1974 2147
rect 2209 2142 2262 2147
rect 2321 2142 2390 2147
rect 2457 2142 2518 2147
rect 2537 2142 2582 2147
rect 2593 2142 2662 2147
rect 2681 2142 2878 2147
rect 2889 2142 2934 2147
rect 961 2137 966 2142
rect 1825 2137 1830 2142
rect 185 2132 270 2137
rect 417 2132 574 2137
rect 569 2127 574 2132
rect 633 2132 758 2137
rect 865 2132 966 2137
rect 1609 2132 1638 2137
rect 1737 2132 1766 2137
rect 1825 2132 2062 2137
rect 2593 2132 2598 2142
rect 2945 2137 2950 2152
rect 3093 2147 3100 2148
rect 3065 2142 3100 2147
rect 3065 2137 3070 2142
rect 3093 2141 3100 2142
rect 2649 2132 2702 2137
rect 2945 2132 3070 2137
rect 633 2127 638 2132
rect 1425 2127 1566 2132
rect 2345 2127 2598 2132
rect 569 2122 638 2127
rect 657 2122 806 2127
rect 825 2122 846 2127
rect 985 2122 1006 2127
rect 1121 2122 1214 2127
rect 1401 2122 1430 2127
rect 1561 2122 2350 2127
rect 2617 2122 2662 2127
rect 2801 2122 2870 2127
rect 801 2117 806 2122
rect 169 2112 214 2117
rect 737 2112 766 2117
rect 801 2112 894 2117
rect 905 2112 974 2117
rect 1113 2112 1198 2117
rect 1217 2112 1294 2117
rect 1385 2112 1414 2117
rect 1409 2107 1414 2112
rect 1473 2112 1550 2117
rect 1473 2107 1478 2112
rect 817 2102 902 2107
rect 993 2102 1158 2107
rect 1273 2102 1334 2107
rect 1409 2102 1478 2107
rect 1497 2102 1526 2107
rect 1545 2097 1550 2112
rect 1777 2112 2030 2117
rect 1777 2097 1782 2112
rect 2025 2107 2030 2112
rect 2361 2112 2798 2117
rect 2361 2107 2366 2112
rect 1801 2102 1846 2107
rect 1945 2102 1982 2107
rect 2025 2102 2366 2107
rect 2385 2102 2510 2107
rect 2625 2102 2734 2107
rect 2889 2102 3006 2107
rect 809 2092 870 2097
rect 977 2092 1006 2097
rect 1089 2092 1118 2097
rect 1545 2092 1782 2097
rect 1833 2092 2006 2097
rect 2801 2092 2942 2097
rect 1001 2087 1094 2092
rect 769 2082 966 2087
rect 961 2077 966 2082
rect 1121 2082 1230 2087
rect 2089 2082 2134 2087
rect 2153 2082 2366 2087
rect 2697 2082 2822 2087
rect 1121 2077 1126 2082
rect 873 2072 902 2077
rect 961 2072 1126 2077
rect 1241 2072 1294 2077
rect 1377 2072 1526 2077
rect 177 2062 198 2067
rect 897 2057 902 2072
rect 1241 2067 1246 2072
rect 1377 2067 1382 2072
rect 1145 2062 1246 2067
rect 1353 2062 1382 2067
rect 1521 2067 1526 2072
rect 1849 2072 2070 2077
rect 1849 2067 1854 2072
rect 1521 2062 1854 2067
rect 2065 2067 2070 2072
rect 2153 2067 2158 2082
rect 2361 2077 2366 2082
rect 2361 2072 2590 2077
rect 2585 2067 2590 2072
rect 2065 2062 2158 2067
rect 2177 2062 2270 2067
rect 2585 2062 2614 2067
rect 1145 2057 1150 2062
rect 1889 2057 2046 2062
rect 2177 2057 2182 2062
rect 897 2052 1150 2057
rect 1417 2052 1502 2057
rect 1865 2052 1894 2057
rect 2041 2052 2182 2057
rect 2265 2057 2270 2062
rect 2265 2052 2934 2057
rect 1417 2047 1422 2052
rect 1497 2047 1846 2052
rect 1169 2042 1422 2047
rect 1841 2042 2254 2047
rect 2745 2042 2766 2047
rect 777 2032 822 2037
rect 1433 2032 1974 2037
rect 2689 2032 2782 2037
rect 2793 2032 2814 2037
rect 2865 2032 2974 2037
rect 2001 2027 2150 2032
rect -7 2017 0 2018
rect 65 2017 70 2027
rect 145 2022 206 2027
rect 425 2022 478 2027
rect 505 2022 542 2027
rect 561 2017 566 2027
rect 665 2022 694 2027
rect 953 2022 1030 2027
rect 1297 2022 1326 2027
rect 1345 2022 1390 2027
rect 1505 2022 1534 2027
rect 1657 2022 1870 2027
rect 1913 2022 1934 2027
rect 1977 2022 2006 2027
rect 2145 2022 2358 2027
rect 2433 2022 2478 2027
rect 2537 2022 2590 2027
rect 2705 2022 2910 2027
rect 3093 2017 3100 2018
rect -7 2012 70 2017
rect 81 2012 110 2017
rect 217 2012 414 2017
rect -7 2011 0 2012
rect 105 2007 222 2012
rect 409 2007 414 2012
rect 545 2012 590 2017
rect 1001 2012 1110 2017
rect 1489 2012 1646 2017
rect 1753 2012 2134 2017
rect 2321 2012 2342 2017
rect 2497 2012 2534 2017
rect 2737 2012 2790 2017
rect 2977 2012 3100 2017
rect 545 2007 550 2012
rect 1641 2007 1758 2012
rect 257 2002 278 2007
rect 409 2002 550 2007
rect 649 2002 758 2007
rect 873 2002 1222 2007
rect 1281 2002 1310 2007
rect 1329 2002 1422 2007
rect 1785 2002 1822 2007
rect 2153 2002 2190 2007
rect 2321 2002 2326 2012
rect 3093 2011 3100 2012
rect 2497 2002 2590 2007
rect 2609 2002 2766 2007
rect -7 1997 0 1998
rect -7 1992 158 1997
rect 849 1992 878 1997
rect 889 1992 926 1997
rect 977 1992 1006 1997
rect 1105 1992 1134 1997
rect -7 1991 0 1992
rect 1001 1987 1110 1992
rect 1217 1987 1222 2002
rect 1329 1997 1334 2002
rect 1241 1992 1334 1997
rect 1417 1997 1422 2002
rect 1913 1997 2086 2002
rect 1417 1992 1446 1997
rect 1457 1992 1518 1997
rect 1537 1992 1646 1997
rect 1705 1992 1766 1997
rect 1777 1992 1798 1997
rect 1889 1992 1918 1997
rect 2081 1992 2110 1997
rect 2265 1992 2342 1997
rect 2417 1992 2462 1997
rect 2545 1992 2646 1997
rect 2777 1992 2798 1997
rect 2809 1992 2846 1997
rect 2865 1992 2918 1997
rect 2161 1987 2246 1992
rect 97 1982 294 1987
rect 313 1982 630 1987
rect 769 1982 886 1987
rect 1217 1982 1614 1987
rect 1745 1982 2062 1987
rect 2121 1982 2166 1987
rect 2241 1982 2446 1987
rect 2489 1982 2790 1987
rect 313 1977 318 1982
rect 185 1972 318 1977
rect 625 1977 630 1982
rect 625 1972 678 1977
rect 817 1972 1662 1977
rect 1745 1967 1750 1982
rect 2057 1977 2126 1982
rect 1769 1972 1798 1977
rect 1833 1972 1870 1977
rect 2177 1972 2278 1977
rect 2337 1972 2390 1977
rect 2401 1972 2430 1977
rect 2689 1972 2766 1977
rect 2849 1972 2894 1977
rect 2425 1967 2566 1972
rect 2689 1967 2694 1972
rect 273 1962 558 1967
rect 585 1962 790 1967
rect 1169 1962 1198 1967
rect 1265 1962 1294 1967
rect 1289 1957 1294 1962
rect 1361 1962 1438 1967
rect 1361 1957 1366 1962
rect 81 1952 190 1957
rect 241 1952 334 1957
rect 497 1952 550 1957
rect 617 1952 686 1957
rect 849 1952 894 1957
rect 929 1952 974 1957
rect 1105 1952 1198 1957
rect 1289 1952 1366 1957
rect 1433 1957 1438 1962
rect 1529 1962 1750 1967
rect 1761 1962 1846 1967
rect 1977 1962 2158 1967
rect 2305 1962 2350 1967
rect 2561 1962 2694 1967
rect 2737 1962 2774 1967
rect 2833 1962 2902 1967
rect 1529 1957 1534 1962
rect 1977 1957 1982 1962
rect 2153 1957 2278 1962
rect 1433 1952 1534 1957
rect 1561 1952 1982 1957
rect 2273 1952 2302 1957
rect 2425 1952 2542 1957
rect 2713 1952 2742 1957
rect 2769 1947 2774 1962
rect 2785 1952 2830 1957
rect 105 1942 206 1947
rect 321 1942 406 1947
rect 433 1942 494 1947
rect 625 1937 630 1947
rect 793 1942 950 1947
rect 961 1942 1014 1947
rect 1161 1942 1190 1947
rect 1385 1942 1414 1947
rect 1553 1942 1630 1947
rect 1729 1942 1838 1947
rect 1881 1942 1918 1947
rect 1993 1942 2070 1947
rect 2089 1942 2134 1947
rect 2161 1942 2294 1947
rect 2313 1942 2374 1947
rect 2441 1942 2478 1947
rect 2537 1942 2638 1947
rect 2705 1942 2734 1947
rect 2769 1942 2830 1947
rect 2913 1942 2958 1947
rect 2289 1937 2294 1942
rect 3093 1937 3100 1938
rect 121 1932 198 1937
rect 217 1932 278 1937
rect 473 1932 534 1937
rect 625 1932 822 1937
rect 833 1932 854 1937
rect 881 1932 942 1937
rect 1073 1932 1118 1937
rect 1169 1932 1862 1937
rect 1921 1932 1990 1937
rect 2145 1932 2182 1937
rect 2289 1932 2326 1937
rect -6 1927 1 1928
rect 817 1927 822 1932
rect 2145 1927 2150 1932
rect 2529 1927 2534 1937
rect 2681 1932 2702 1937
rect 3009 1932 3100 1937
rect 3093 1931 3100 1932
rect -6 1922 134 1927
rect 289 1922 454 1927
rect 521 1922 670 1927
rect 817 1922 1030 1927
rect 1057 1922 1182 1927
rect 1353 1922 1478 1927
rect 1593 1922 1662 1927
rect 1745 1922 1774 1927
rect 1913 1922 1998 1927
rect 2129 1922 2150 1927
rect 2409 1922 2454 1927
rect 2497 1922 2534 1927
rect 2673 1922 2750 1927
rect 2913 1922 2998 1927
rect -6 1921 1 1922
rect 129 1912 134 1922
rect 3093 1917 3100 1918
rect 201 1912 318 1917
rect 329 1912 438 1917
rect 513 1912 614 1917
rect 641 1912 702 1917
rect 857 1912 886 1917
rect 969 1912 1062 1917
rect 1105 1912 1262 1917
rect 1433 1912 1510 1917
rect 1793 1912 2006 1917
rect 2161 1912 2190 1917
rect 2321 1912 2446 1917
rect 2537 1912 2582 1917
rect 2713 1912 2798 1917
rect 3025 1912 3100 1917
rect -6 1907 1 1908
rect 1105 1907 1110 1912
rect 1705 1907 1774 1912
rect 3093 1911 3100 1912
rect -6 1902 86 1907
rect 425 1902 478 1907
rect 529 1902 598 1907
rect 625 1902 1110 1907
rect 1121 1902 1182 1907
rect 1233 1902 1278 1907
rect 1617 1902 1710 1907
rect 1769 1902 2174 1907
rect 2713 1902 2742 1907
rect 2873 1902 2934 1907
rect -6 1901 1 1902
rect 593 1897 598 1902
rect 217 1892 286 1897
rect 465 1892 582 1897
rect 593 1892 694 1897
rect 977 1892 1246 1897
rect 1297 1892 1374 1897
rect 1721 1892 1838 1897
rect 1297 1887 1302 1892
rect 289 1882 478 1887
rect 473 1877 478 1882
rect 777 1882 934 1887
rect 953 1882 1022 1887
rect 1081 1882 1126 1887
rect 1153 1882 1182 1887
rect 1249 1882 1302 1887
rect 1369 1887 1374 1892
rect 1833 1887 1838 1892
rect 1929 1892 2006 1897
rect 2129 1892 2158 1897
rect 1929 1887 1934 1892
rect 2001 1887 2134 1892
rect 2737 1887 2806 1892
rect 1369 1882 1398 1887
rect 1601 1882 1710 1887
rect 1833 1882 1934 1887
rect 1953 1882 1982 1887
rect 2281 1882 2302 1887
rect 2521 1882 2742 1887
rect 2801 1882 2862 1887
rect 777 1877 782 1882
rect 473 1872 678 1877
rect 689 1872 782 1877
rect 929 1877 934 1882
rect 1705 1877 1814 1882
rect 929 1872 1214 1877
rect 1369 1872 1446 1877
rect 345 1862 454 1867
rect 345 1857 350 1862
rect 321 1852 350 1857
rect 449 1857 454 1862
rect 673 1857 678 1872
rect 1809 1867 1814 1877
rect 1953 1867 1958 1882
rect 2857 1877 2862 1882
rect 2945 1882 3030 1887
rect 2945 1877 2950 1882
rect 2089 1872 2198 1877
rect 2753 1872 2790 1877
rect 2857 1872 2950 1877
rect 793 1862 1014 1867
rect 793 1857 798 1862
rect 1009 1857 1014 1862
rect 1097 1862 1150 1867
rect 1209 1862 1398 1867
rect 1097 1857 1102 1862
rect 449 1852 630 1857
rect 673 1852 798 1857
rect 865 1852 990 1857
rect 1009 1852 1102 1857
rect 1393 1857 1398 1862
rect 1457 1862 1718 1867
rect 1809 1862 1958 1867
rect 2049 1862 2310 1867
rect 1457 1857 1462 1862
rect 1393 1852 1462 1857
rect 2681 1852 2710 1857
rect 345 1842 486 1847
rect 1121 1842 1166 1847
rect 1689 1842 1790 1847
rect 2081 1842 2182 1847
rect 2081 1837 2086 1842
rect 305 1832 326 1837
rect 393 1832 422 1837
rect 505 1832 534 1837
rect 817 1832 894 1837
rect 1009 1832 1118 1837
rect 1145 1832 1430 1837
rect 1497 1832 1766 1837
rect 1857 1832 1886 1837
rect 2057 1832 2086 1837
rect 2177 1837 2182 1842
rect 2393 1842 2470 1847
rect 2809 1842 2862 1847
rect 2393 1837 2398 1842
rect 2177 1832 2342 1837
rect 2369 1832 2398 1837
rect 2465 1837 2470 1842
rect 2465 1832 2518 1837
rect 2617 1832 2694 1837
rect 2849 1832 2918 1837
rect 89 1822 126 1827
rect 409 1822 446 1827
rect 353 1812 430 1817
rect 465 1807 470 1827
rect 737 1822 870 1827
rect 993 1822 1054 1827
rect 1297 1822 1334 1827
rect 1433 1822 1574 1827
rect 1745 1822 1886 1827
rect 2025 1822 2070 1827
rect 2121 1822 2214 1827
rect 2321 1822 2350 1827
rect 2409 1822 2486 1827
rect 2761 1822 2814 1827
rect 2345 1817 2414 1822
rect 497 1812 590 1817
rect 785 1812 814 1817
rect 881 1812 1102 1817
rect 1129 1812 1166 1817
rect 1201 1812 1254 1817
rect 1265 1812 1358 1817
rect 1449 1812 1486 1817
rect 1561 1812 1702 1817
rect 1737 1812 1950 1817
rect 2009 1812 2070 1817
rect 2089 1812 2118 1817
rect 2745 1812 2782 1817
rect 809 1807 886 1812
rect 1697 1807 1702 1812
rect 97 1802 182 1807
rect 417 1802 470 1807
rect 585 1802 654 1807
rect 961 1802 1006 1807
rect 1129 1802 1230 1807
rect 1697 1802 2054 1807
rect 2065 1802 2070 1812
rect 2305 1802 2334 1807
rect 2345 1802 2518 1807
rect 1249 1797 1358 1802
rect 137 1792 166 1797
rect 297 1792 422 1797
rect 441 1792 494 1797
rect 641 1792 702 1797
rect 833 1792 998 1797
rect 1097 1792 1254 1797
rect 1353 1792 1518 1797
rect 1529 1792 1726 1797
rect 1753 1792 1814 1797
rect 1825 1792 1894 1797
rect 1953 1792 2030 1797
rect 2313 1792 2414 1797
rect 2657 1792 2702 1797
rect 2833 1792 2878 1797
rect 417 1787 422 1792
rect 145 1782 246 1787
rect 417 1782 502 1787
rect 537 1782 678 1787
rect 697 1782 774 1787
rect 913 1782 934 1787
rect 1225 1782 1342 1787
rect 1713 1782 2062 1787
rect 2209 1782 2302 1787
rect 2297 1777 2302 1782
rect 2361 1782 2390 1787
rect 2801 1782 2878 1787
rect 2361 1777 2366 1782
rect 265 1772 358 1777
rect 793 1772 822 1777
rect 1193 1772 1374 1777
rect 1769 1772 1958 1777
rect 2017 1772 2046 1777
rect 2297 1772 2366 1777
rect 265 1767 270 1772
rect 81 1762 150 1767
rect 193 1762 270 1767
rect 353 1767 358 1772
rect 425 1767 614 1772
rect 857 1767 942 1772
rect 1953 1767 1958 1772
rect 353 1762 430 1767
rect 609 1762 862 1767
rect 937 1762 1070 1767
rect 1273 1762 1294 1767
rect 1569 1762 1670 1767
rect 1857 1762 1934 1767
rect 1953 1762 2126 1767
rect 2153 1762 2230 1767
rect 2385 1762 2558 1767
rect 2769 1762 2822 1767
rect 145 1757 150 1762
rect 2153 1757 2158 1762
rect 73 1752 126 1757
rect 145 1752 342 1757
rect 337 1747 342 1752
rect 441 1752 542 1757
rect 561 1752 630 1757
rect 873 1752 926 1757
rect 1265 1752 1326 1757
rect 1465 1752 1510 1757
rect 1745 1752 2158 1757
rect 2225 1757 2230 1762
rect 2225 1752 2302 1757
rect 441 1747 446 1752
rect 113 1742 318 1747
rect 337 1742 446 1747
rect 489 1742 590 1747
rect 617 1742 782 1747
rect 817 1742 846 1747
rect 969 1742 1078 1747
rect 1257 1742 1286 1747
rect 1657 1742 1702 1747
rect 1865 1742 1894 1747
rect 1905 1742 2094 1747
rect 2169 1742 2214 1747
rect 2329 1742 2462 1747
rect 2553 1742 2598 1747
rect 2785 1742 2814 1747
rect 2865 1742 2950 1747
rect 169 1732 246 1737
rect 265 1732 302 1737
rect 465 1732 814 1737
rect 1025 1732 1142 1737
rect 1169 1732 1206 1737
rect 1361 1732 1398 1737
rect 1721 1732 1774 1737
rect 1361 1727 1366 1732
rect 1889 1727 1894 1742
rect 2193 1727 2198 1737
rect 2353 1732 2414 1737
rect 2465 1732 2494 1737
rect 2913 1732 3014 1737
rect 217 1722 262 1727
rect 305 1722 358 1727
rect 481 1722 534 1727
rect 625 1722 654 1727
rect 729 1722 806 1727
rect 841 1722 886 1727
rect 529 1717 630 1722
rect 913 1717 918 1727
rect 1073 1722 1190 1727
rect 1281 1722 1366 1727
rect 1377 1722 1414 1727
rect 1585 1722 1694 1727
rect 1889 1722 1910 1727
rect 2049 1722 2094 1727
rect 2169 1722 2198 1727
rect 2257 1722 2358 1727
rect 2857 1722 2886 1727
rect 1073 1717 1078 1722
rect 2897 1717 2902 1727
rect 65 1712 510 1717
rect 681 1712 726 1717
rect 833 1712 918 1717
rect 1017 1712 1078 1717
rect 1209 1712 1262 1717
rect 1297 1712 1350 1717
rect 1641 1712 1670 1717
rect 1705 1712 1990 1717
rect 2249 1712 2278 1717
rect 2273 1707 2278 1712
rect 2401 1712 2494 1717
rect 2585 1712 2630 1717
rect 2897 1712 2918 1717
rect 2401 1707 2406 1712
rect 353 1702 478 1707
rect 553 1702 662 1707
rect 705 1702 742 1707
rect 769 1702 918 1707
rect 1089 1702 1238 1707
rect 1305 1702 1366 1707
rect 1561 1702 1702 1707
rect 1897 1702 1958 1707
rect 2273 1702 2406 1707
rect 2609 1702 2630 1707
rect 2857 1702 2902 1707
rect 553 1697 558 1702
rect 505 1692 558 1697
rect 657 1697 662 1702
rect 657 1692 1046 1697
rect 1185 1692 1278 1697
rect 1425 1692 1510 1697
rect 1881 1692 1926 1697
rect 2905 1692 2958 1697
rect 1425 1687 1430 1692
rect 569 1682 1126 1687
rect 1249 1682 1278 1687
rect 1273 1677 1278 1682
rect 1377 1682 1430 1687
rect 1505 1687 1510 1692
rect 1505 1682 1534 1687
rect 1873 1682 1910 1687
rect 2425 1682 2446 1687
rect 2505 1682 2566 1687
rect 1377 1677 1382 1682
rect 457 1672 998 1677
rect 1049 1672 1086 1677
rect 1273 1672 1382 1677
rect 1441 1672 1470 1677
rect 1465 1667 1470 1672
rect 1545 1672 1862 1677
rect 1921 1672 2230 1677
rect 1545 1667 1550 1672
rect 1857 1667 1926 1672
rect 553 1662 598 1667
rect 593 1657 598 1662
rect 689 1662 1094 1667
rect 1465 1662 1550 1667
rect 689 1657 694 1662
rect 305 1652 406 1657
rect 593 1652 694 1657
rect 713 1652 742 1657
rect 881 1652 1150 1657
rect 1817 1652 1942 1657
rect 2753 1652 2870 1657
rect 2889 1652 2958 1657
rect 305 1647 310 1652
rect 241 1642 310 1647
rect 401 1647 406 1652
rect 737 1647 886 1652
rect 2889 1647 2894 1652
rect 401 1642 574 1647
rect 905 1642 958 1647
rect 1009 1642 1182 1647
rect 1321 1642 1366 1647
rect 1569 1642 1654 1647
rect 2225 1642 2318 1647
rect 2665 1642 2806 1647
rect 2841 1642 2894 1647
rect 2953 1647 2958 1652
rect 2953 1642 2982 1647
rect 2225 1637 2230 1642
rect 257 1632 390 1637
rect 681 1632 798 1637
rect 897 1632 942 1637
rect 1105 1632 1142 1637
rect 1265 1632 1334 1637
rect 1345 1632 1390 1637
rect 1417 1632 1550 1637
rect 1561 1632 1598 1637
rect 1697 1632 1806 1637
rect 1345 1627 1350 1632
rect 1801 1627 1806 1632
rect 1889 1632 2230 1637
rect 2313 1637 2318 1642
rect 2313 1632 2382 1637
rect 2625 1632 2750 1637
rect 2761 1632 2790 1637
rect 2849 1632 2878 1637
rect 1889 1627 1894 1632
rect 177 1622 326 1627
rect 537 1622 606 1627
rect 825 1622 918 1627
rect 1073 1622 1142 1627
rect 1297 1622 1350 1627
rect 1377 1622 1462 1627
rect 1537 1622 1574 1627
rect 1633 1622 1662 1627
rect 1801 1622 1894 1627
rect 1913 1622 1998 1627
rect 2025 1622 2062 1627
rect 2209 1622 2278 1627
rect 2297 1622 2326 1627
rect 2369 1622 2430 1627
rect 2585 1622 2638 1627
rect 2793 1622 2830 1627
rect 2913 1622 3014 1627
rect 2081 1617 2190 1622
rect 145 1612 190 1617
rect 409 1612 478 1617
rect 729 1612 758 1617
rect 1257 1612 1390 1617
rect 1401 1612 1470 1617
rect 1577 1612 1606 1617
rect 1985 1612 2086 1617
rect 2185 1612 2254 1617
rect 2385 1612 2478 1617
rect 2721 1612 2742 1617
rect 2785 1612 2830 1617
rect 409 1607 414 1612
rect 161 1602 182 1607
rect 225 1602 414 1607
rect 473 1607 478 1612
rect 473 1602 558 1607
rect 577 1602 630 1607
rect 713 1602 750 1607
rect 1129 1602 1158 1607
rect 1417 1602 1446 1607
rect 1625 1602 1742 1607
rect 2041 1602 2206 1607
rect 2289 1602 2366 1607
rect 2513 1602 2646 1607
rect 81 1592 110 1597
rect 129 1592 190 1597
rect 209 1592 302 1597
rect 313 1592 390 1597
rect 433 1592 462 1597
rect 577 1592 582 1602
rect 2201 1597 2294 1602
rect 633 1592 806 1597
rect 1609 1592 1638 1597
rect 1713 1592 1950 1597
rect 2697 1592 2742 1597
rect 2785 1592 2854 1597
rect 81 1582 126 1587
rect 697 1582 886 1587
rect 1161 1582 1334 1587
rect 1513 1582 1622 1587
rect 2161 1582 2190 1587
rect 2369 1582 2438 1587
rect 2505 1582 2686 1587
rect 2865 1582 2934 1587
rect 2681 1577 2870 1582
rect 673 1572 790 1577
rect 785 1567 790 1572
rect 873 1572 902 1577
rect 1185 1572 1262 1577
rect 1617 1572 1654 1577
rect 2041 1572 2102 1577
rect 2249 1572 2406 1577
rect 873 1567 878 1572
rect 1281 1567 1414 1572
rect 361 1562 398 1567
rect 785 1562 878 1567
rect 1241 1562 1286 1567
rect 1409 1562 1438 1567
rect 1529 1562 1630 1567
rect 1641 1562 1774 1567
rect 1937 1562 2022 1567
rect 2089 1562 2294 1567
rect 2577 1562 2726 1567
rect 2753 1562 2838 1567
rect 2881 1562 2934 1567
rect 273 1552 470 1557
rect 609 1552 766 1557
rect 1129 1552 1294 1557
rect 1305 1552 1374 1557
rect 1665 1552 1694 1557
rect 1937 1552 2118 1557
rect 2209 1552 2262 1557
rect 2409 1552 2502 1557
rect 2705 1552 2854 1557
rect 2113 1547 2118 1552
rect 129 1542 206 1547
rect 241 1527 246 1547
rect 281 1542 366 1547
rect 561 1542 622 1547
rect 297 1532 318 1537
rect 337 1532 390 1537
rect 705 1527 710 1547
rect 793 1542 854 1547
rect 929 1542 990 1547
rect 1193 1542 1390 1547
rect 1601 1542 1662 1547
rect 1761 1542 1806 1547
rect 1905 1542 1974 1547
rect 1993 1542 2094 1547
rect 2113 1542 2222 1547
rect 2249 1542 2318 1547
rect 2425 1542 2502 1547
rect 2641 1542 2742 1547
rect 2833 1542 2902 1547
rect 1969 1537 1974 1542
rect 1225 1532 1254 1537
rect 1361 1532 1398 1537
rect 1905 1532 1942 1537
rect 1969 1532 2198 1537
rect 2697 1532 2774 1537
rect 217 1522 246 1527
rect 513 1522 606 1527
rect 705 1522 790 1527
rect 841 1522 878 1527
rect 1305 1522 1358 1527
rect 353 1512 422 1517
rect 561 1512 646 1517
rect 761 1512 942 1517
rect 1201 1512 1310 1517
rect 1321 1512 1390 1517
rect 1473 1507 1478 1527
rect 1681 1522 1766 1527
rect 1585 1512 1614 1517
rect 1905 1512 1910 1532
rect 1977 1522 2006 1527
rect 2161 1522 2254 1527
rect 2337 1522 2382 1527
rect 2401 1522 2454 1527
rect 2777 1522 2814 1527
rect 2001 1517 2166 1522
rect 1937 1512 1966 1517
rect 2185 1512 2214 1517
rect 2273 1512 2374 1517
rect 2385 1512 2462 1517
rect 2545 1512 2798 1517
rect 2889 1512 2918 1517
rect 2545 1507 2550 1512
rect 857 1502 934 1507
rect 1265 1502 1326 1507
rect 1473 1502 1606 1507
rect 1785 1502 1854 1507
rect 1969 1502 2238 1507
rect 1785 1497 1790 1502
rect 769 1492 1030 1497
rect 1369 1492 1430 1497
rect 1545 1492 1790 1497
rect 1849 1497 1854 1502
rect 2233 1497 2238 1502
rect 2345 1502 2550 1507
rect 2801 1502 2870 1507
rect 2345 1497 2350 1502
rect 1849 1492 1894 1497
rect 1889 1487 1894 1492
rect 2129 1492 2206 1497
rect 2233 1492 2350 1497
rect 2369 1492 2446 1497
rect 2849 1492 2894 1497
rect 1521 1482 1550 1487
rect 1545 1477 1550 1482
rect 1673 1482 1702 1487
rect 1777 1482 1838 1487
rect 1889 1482 1958 1487
rect 1673 1477 1678 1482
rect 1545 1472 1678 1477
rect 1953 1477 1958 1482
rect 2129 1477 2134 1492
rect 2153 1482 2214 1487
rect 2561 1482 2606 1487
rect 2761 1482 2798 1487
rect 1953 1472 2134 1477
rect 2449 1472 2638 1477
rect 2689 1472 2766 1477
rect 2881 1472 2966 1477
rect 1257 1462 1334 1467
rect 1257 1457 1262 1462
rect 665 1452 702 1457
rect 1185 1452 1262 1457
rect 1329 1457 1334 1462
rect 2233 1462 2430 1467
rect 1329 1452 1486 1457
rect 1713 1452 1870 1457
rect 2233 1447 2238 1462
rect 2425 1457 2430 1462
rect 2425 1452 2534 1457
rect 713 1442 950 1447
rect 1953 1442 2038 1447
rect 2201 1442 2238 1447
rect 2529 1447 2534 1452
rect 2529 1442 2758 1447
rect 329 1432 478 1437
rect 769 1432 1006 1437
rect 1273 1432 1318 1437
rect 1433 1432 1478 1437
rect 1953 1432 1982 1437
rect 1977 1427 1982 1432
rect 2049 1432 2078 1437
rect 2113 1432 2190 1437
rect 2049 1427 2054 1432
rect 2185 1427 2190 1432
rect 2249 1432 2318 1437
rect 2417 1432 2518 1437
rect 2777 1432 2902 1437
rect 2249 1427 2254 1432
rect 2777 1427 2782 1432
rect 161 1422 198 1427
rect 809 1422 846 1427
rect 929 1422 966 1427
rect 1057 1422 1166 1427
rect 1201 1422 1238 1427
rect 1321 1422 1342 1427
rect 1977 1422 2054 1427
rect 2097 1422 2134 1427
rect 2185 1422 2254 1427
rect 2489 1422 2542 1427
rect 2601 1422 2782 1427
rect 2897 1427 2902 1432
rect 2897 1422 2926 1427
rect 1057 1417 1062 1422
rect 225 1412 294 1417
rect 369 1412 430 1417
rect 593 1412 678 1417
rect 985 1412 1062 1417
rect 1297 1412 1358 1417
rect 2081 1412 2126 1417
rect 2289 1412 2366 1417
rect 2401 1412 2462 1417
rect 2553 1412 2598 1417
rect 2609 1412 2630 1417
rect 2697 1412 2958 1417
rect 593 1407 598 1412
rect 305 1402 326 1407
rect 569 1402 598 1407
rect 673 1407 678 1412
rect 673 1402 702 1407
rect 761 1402 790 1407
rect 993 1402 1022 1407
rect 1017 1397 1022 1402
rect 1169 1402 1206 1407
rect 1297 1402 1350 1407
rect 1617 1402 1654 1407
rect 1865 1402 1894 1407
rect 2113 1402 2270 1407
rect 1169 1397 1174 1402
rect 2289 1397 2294 1412
rect 2361 1407 2366 1412
rect 2361 1402 2654 1407
rect 289 1392 350 1397
rect 425 1392 646 1397
rect 689 1392 726 1397
rect 801 1392 886 1397
rect 1017 1392 1174 1397
rect 1193 1392 1374 1397
rect 1497 1392 1558 1397
rect 1697 1392 1814 1397
rect 1953 1392 1998 1397
rect 2065 1392 2110 1397
rect 2209 1392 2294 1397
rect 2305 1392 2350 1397
rect 2425 1392 2590 1397
rect 2753 1392 2774 1397
rect 641 1387 646 1392
rect 321 1382 358 1387
rect 641 1382 790 1387
rect 785 1377 790 1382
rect 897 1382 990 1387
rect 1337 1382 1398 1387
rect 1793 1382 1822 1387
rect 897 1377 902 1382
rect 1817 1377 1822 1382
rect 1913 1382 1950 1387
rect 2169 1382 2222 1387
rect 2273 1382 2318 1387
rect 2393 1382 2702 1387
rect 1913 1377 1918 1382
rect 2785 1377 2790 1407
rect 2833 1382 2974 1387
rect 225 1372 318 1377
rect 785 1372 902 1377
rect 1201 1372 1230 1377
rect 1225 1367 1230 1372
rect 1337 1372 1366 1377
rect 1817 1372 1918 1377
rect 2137 1372 2334 1377
rect 2425 1372 2526 1377
rect 2577 1372 2742 1377
rect 2769 1372 2790 1377
rect 1337 1367 1342 1372
rect 137 1362 206 1367
rect 1049 1362 1094 1367
rect 1169 1362 1206 1367
rect 1225 1362 1342 1367
rect 1545 1362 1734 1367
rect 1937 1362 1966 1367
rect 2137 1362 2358 1367
rect 2385 1362 2494 1367
rect 2513 1362 2542 1367
rect 2609 1362 2742 1367
rect 2833 1362 2878 1367
rect 2385 1357 2390 1362
rect 161 1352 182 1357
rect 585 1352 998 1357
rect 1033 1352 1174 1357
rect 1497 1352 1518 1357
rect 1561 1352 1590 1357
rect 1713 1352 1758 1357
rect 2017 1352 2070 1357
rect 2225 1352 2390 1357
rect 2401 1352 2630 1357
rect 2657 1352 2806 1357
rect 153 1342 390 1347
rect 601 1342 654 1347
rect 1025 1342 1070 1347
rect 1361 1342 1494 1347
rect 1513 1342 1574 1347
rect 1665 1342 1718 1347
rect 1881 1342 2006 1347
rect 2049 1342 2110 1347
rect 2433 1342 2518 1347
rect 209 1332 262 1337
rect 561 1332 630 1337
rect 857 1332 902 1337
rect 1009 1332 1078 1337
rect 89 1322 326 1327
rect 409 1322 430 1327
rect 473 1322 510 1327
rect 529 1322 566 1327
rect 601 1322 638 1327
rect 1289 1322 1446 1327
rect 1481 1322 1518 1327
rect 1681 1322 1686 1342
rect 2337 1332 2454 1337
rect 1937 1327 2102 1332
rect 2561 1327 2566 1347
rect 2585 1342 2686 1347
rect 2705 1342 2750 1347
rect 2849 1342 2998 1347
rect 2601 1332 2638 1337
rect 2673 1327 2678 1337
rect 2713 1332 2878 1337
rect 1849 1322 1942 1327
rect 2097 1322 2126 1327
rect 2561 1322 2654 1327
rect 2673 1322 2694 1327
rect 2729 1322 2822 1327
rect 81 1312 110 1317
rect 209 1312 238 1317
rect 321 1312 326 1322
rect 337 1312 374 1317
rect 497 1312 542 1317
rect 561 1312 566 1322
rect 713 1312 750 1317
rect 921 1312 966 1317
rect 1321 1312 1358 1317
rect 1489 1312 1646 1317
rect 1777 1312 1846 1317
rect 1929 1312 1982 1317
rect 2041 1312 2086 1317
rect 2457 1312 2606 1317
rect 2625 1312 2678 1317
rect 2769 1312 2854 1317
rect 2905 1312 2934 1317
rect 105 1307 214 1312
rect 249 1302 270 1307
rect 401 1302 486 1307
rect 857 1302 902 1307
rect 1225 1302 1278 1307
rect 1273 1297 1278 1302
rect 1401 1302 1478 1307
rect 1713 1302 1766 1307
rect 1401 1297 1406 1302
rect 1761 1297 1766 1302
rect 1833 1302 1886 1307
rect 1833 1297 1838 1302
rect 177 1292 302 1297
rect 313 1292 454 1297
rect 465 1292 558 1297
rect 1009 1292 1118 1297
rect 1273 1292 1406 1297
rect 1457 1292 1526 1297
rect 1761 1292 1838 1297
rect 1881 1297 1886 1302
rect 1953 1302 2166 1307
rect 2273 1302 2438 1307
rect 2473 1302 2502 1307
rect 1953 1297 1958 1302
rect 2497 1297 2502 1302
rect 2593 1302 2718 1307
rect 2745 1302 2790 1307
rect 2593 1297 2598 1302
rect 1881 1292 1958 1297
rect 2001 1292 2046 1297
rect 2249 1292 2278 1297
rect 2497 1292 2598 1297
rect 2617 1292 2782 1297
rect 2809 1292 2926 1297
rect 449 1287 454 1292
rect 273 1282 334 1287
rect 449 1282 598 1287
rect 1425 1282 1454 1287
rect 329 1277 438 1282
rect 1449 1277 1454 1282
rect 1521 1282 1550 1287
rect 2281 1282 2318 1287
rect 1521 1277 1526 1282
rect 233 1272 310 1277
rect 433 1272 582 1277
rect 1449 1272 1526 1277
rect 2065 1272 2230 1277
rect 2065 1267 2070 1272
rect 161 1262 494 1267
rect 609 1262 710 1267
rect 1985 1262 2070 1267
rect 2225 1267 2230 1272
rect 2417 1272 2598 1277
rect 2777 1272 2894 1277
rect 2417 1267 2422 1272
rect 2225 1262 2358 1267
rect 2393 1262 2422 1267
rect 2593 1267 2598 1272
rect 2593 1262 2686 1267
rect 169 1252 222 1257
rect 297 1252 334 1257
rect 409 1252 486 1257
rect 2089 1252 2206 1257
rect 2345 1252 2398 1257
rect 2441 1252 2462 1257
rect 2489 1252 2526 1257
rect 2569 1252 2622 1257
rect 2705 1252 2742 1257
rect 2089 1247 2094 1252
rect 97 1242 182 1247
rect 217 1242 326 1247
rect 345 1242 422 1247
rect 817 1242 990 1247
rect 1009 1242 1086 1247
rect 1009 1237 1014 1242
rect 121 1232 198 1237
rect 273 1232 382 1237
rect 449 1232 478 1237
rect 697 1232 870 1237
rect 977 1232 1014 1237
rect 1081 1237 1086 1242
rect 1873 1242 1966 1247
rect 2033 1242 2094 1247
rect 2201 1247 2206 1252
rect 2201 1242 2230 1247
rect 1873 1237 1878 1242
rect 1081 1232 1110 1237
rect 1161 1232 1502 1237
rect 1601 1232 1678 1237
rect 1849 1232 1878 1237
rect 1961 1237 1966 1242
rect 1961 1232 2118 1237
rect 2169 1232 2286 1237
rect 2313 1232 2334 1237
rect 2361 1232 2478 1237
rect 2545 1232 2614 1237
rect 2769 1232 2790 1237
rect 2545 1227 2550 1232
rect 129 1222 190 1227
rect 209 1217 214 1227
rect 281 1222 318 1227
rect 353 1222 534 1227
rect 665 1222 742 1227
rect 817 1222 886 1227
rect 969 1222 1038 1227
rect 1081 1222 1134 1227
rect 1153 1222 1198 1227
rect 1265 1222 1286 1227
rect 1825 1222 1902 1227
rect 1969 1222 1990 1227
rect 2089 1222 2150 1227
rect 2497 1222 2550 1227
rect 2593 1222 2630 1227
rect 2737 1222 2766 1227
rect 185 1212 214 1217
rect 241 1212 358 1217
rect 393 1212 438 1217
rect 489 1212 518 1217
rect 1833 1212 1870 1217
rect 1905 1212 1926 1217
rect 2641 1212 2678 1217
rect 2713 1212 2758 1217
rect 2785 1212 2822 1217
rect 241 1202 270 1207
rect 265 1197 270 1202
rect 369 1202 446 1207
rect 1273 1202 1398 1207
rect 1569 1202 1598 1207
rect 1649 1202 1726 1207
rect 1921 1202 1926 1212
rect 2065 1202 2158 1207
rect 2681 1202 2838 1207
rect 369 1197 374 1202
rect 265 1192 374 1197
rect 393 1192 422 1197
rect 417 1187 422 1192
rect 529 1192 646 1197
rect 689 1192 742 1197
rect 761 1192 838 1197
rect 857 1192 926 1197
rect 1217 1192 1310 1197
rect 1385 1192 1454 1197
rect 1625 1192 1694 1197
rect 1825 1192 1894 1197
rect 1913 1192 1934 1197
rect 1953 1192 2150 1197
rect 2169 1192 2214 1197
rect 2385 1192 2422 1197
rect 2473 1192 2542 1197
rect 2593 1192 2758 1197
rect 2905 1192 2950 1197
rect 529 1187 534 1192
rect 417 1182 534 1187
rect 737 1187 742 1192
rect 1953 1187 1958 1192
rect 737 1182 1014 1187
rect 1073 1182 1134 1187
rect 1249 1182 1286 1187
rect 1521 1182 1646 1187
rect 1641 1177 1646 1182
rect 1737 1182 1814 1187
rect 1905 1182 1958 1187
rect 2025 1182 2166 1187
rect 2225 1182 2302 1187
rect 2449 1182 2534 1187
rect 2697 1182 2822 1187
rect 1737 1177 1742 1182
rect 2161 1177 2230 1182
rect 633 1172 726 1177
rect 753 1172 822 1177
rect 873 1172 998 1177
rect 1201 1172 1446 1177
rect 1529 1172 1590 1177
rect 1641 1172 1742 1177
rect 2105 1172 2142 1177
rect 2417 1172 2558 1177
rect 2617 1172 2702 1177
rect 2873 1172 2918 1177
rect 193 1162 262 1167
rect 721 1162 1174 1167
rect 1289 1162 1326 1167
rect 1801 1162 1838 1167
rect 2009 1162 2182 1167
rect 2441 1162 2630 1167
rect 2721 1162 2838 1167
rect 601 1157 694 1162
rect 2625 1157 2726 1162
rect 2833 1157 2838 1162
rect 161 1152 182 1157
rect 409 1152 550 1157
rect 577 1152 606 1157
rect 689 1152 846 1157
rect 841 1147 846 1152
rect 985 1152 1054 1157
rect 1441 1152 1622 1157
rect 1873 1152 2102 1157
rect 2545 1152 2606 1157
rect 2833 1152 2894 1157
rect 985 1147 990 1152
rect 177 1142 286 1147
rect 393 1142 454 1147
rect 545 1142 678 1147
rect 745 1142 822 1147
rect 841 1142 990 1147
rect 1009 1142 1094 1147
rect 1401 1142 1486 1147
rect 1577 1142 1694 1147
rect 1993 1142 2030 1147
rect 2057 1142 2118 1147
rect 2161 1142 2206 1147
rect 2337 1142 2438 1147
rect 2513 1142 2582 1147
rect 2625 1142 2662 1147
rect 2769 1142 2806 1147
rect 2881 1142 2926 1147
rect 369 1132 470 1137
rect 537 1132 630 1137
rect 657 1132 750 1137
rect 1825 1132 1886 1137
rect 2585 1132 2646 1137
rect 2785 1132 2830 1137
rect 209 1122 342 1127
rect 601 1122 726 1127
rect 1065 1122 1118 1127
rect 1465 1122 1494 1127
rect 1889 1122 2134 1127
rect 2305 1122 2454 1127
rect 2537 1122 2598 1127
rect 2625 1122 2774 1127
rect 2857 1122 2950 1127
rect 2593 1117 2598 1122
rect 305 1112 390 1117
rect 409 1112 526 1117
rect 545 1112 662 1117
rect 825 1112 934 1117
rect 993 1112 1054 1117
rect 1217 1112 1262 1117
rect 1473 1112 1558 1117
rect 1897 1112 1934 1117
rect 2137 1112 2182 1117
rect 2257 1112 2326 1117
rect 2473 1112 2502 1117
rect 2593 1112 2646 1117
rect 2665 1112 2726 1117
rect 2865 1112 2894 1117
rect 297 1102 350 1107
rect 497 1102 542 1107
rect 609 1102 878 1107
rect 1329 1102 1470 1107
rect 1545 1102 1622 1107
rect 2161 1102 2270 1107
rect 2297 1102 2358 1107
rect 2353 1097 2358 1102
rect 2489 1102 2518 1107
rect 2697 1102 2782 1107
rect 2817 1102 2926 1107
rect 2489 1097 2494 1102
rect 625 1092 654 1097
rect 417 1082 518 1087
rect 649 1077 654 1092
rect 841 1092 910 1097
rect 1073 1092 1206 1097
rect 841 1077 846 1092
rect 1201 1087 1206 1092
rect 1273 1092 1318 1097
rect 1273 1087 1278 1092
rect 929 1082 998 1087
rect 1201 1082 1278 1087
rect 1313 1087 1318 1092
rect 1377 1092 1406 1097
rect 1961 1092 2286 1097
rect 2305 1092 2334 1097
rect 2353 1092 2494 1097
rect 2833 1092 2926 1097
rect 1377 1087 1382 1092
rect 1313 1082 1382 1087
rect 1641 1082 1886 1087
rect 2225 1082 2286 1087
rect 929 1077 934 1082
rect 649 1072 846 1077
rect 865 1072 934 1077
rect 993 1077 998 1082
rect 993 1072 1022 1077
rect 1641 1067 1646 1082
rect 929 1062 1054 1067
rect 1593 1062 1646 1067
rect 1881 1067 1886 1082
rect 2601 1072 2622 1077
rect 2865 1072 2982 1077
rect 1881 1062 2110 1067
rect 921 1052 982 1057
rect 1649 1052 1870 1057
rect 2169 1052 2222 1057
rect 2345 1052 2486 1057
rect 289 1042 382 1047
rect 897 1042 982 1047
rect 1049 1042 1142 1047
rect 1633 1042 1694 1047
rect 2625 1042 2710 1047
rect 161 1032 206 1037
rect 369 1032 462 1037
rect 529 1032 566 1037
rect 841 1032 894 1037
rect 1033 1032 1102 1037
rect 1673 1032 1734 1037
rect 1921 1032 2006 1037
rect 2193 1032 2310 1037
rect 2337 1032 2366 1037
rect 2641 1032 2678 1037
rect 2689 1032 2718 1037
rect 2761 1032 2790 1037
rect 137 1022 182 1027
rect 209 1022 254 1027
rect 337 1022 430 1027
rect 665 1022 766 1027
rect 873 1022 1062 1027
rect 1201 1022 1270 1027
rect 1289 1022 1318 1027
rect 1337 1022 1390 1027
rect 1473 1022 1502 1027
rect 1609 1022 1742 1027
rect 1921 1022 2030 1027
rect 2041 1022 2150 1027
rect 2505 1022 2606 1027
rect 121 1012 166 1017
rect 417 1012 582 1017
rect 849 1012 902 1017
rect 985 1012 1206 1017
rect 1249 1012 1430 1017
rect 1585 1012 1686 1017
rect 1905 1012 2038 1017
rect 2065 1012 2086 1017
rect 2417 1012 2478 1017
rect 745 1007 822 1012
rect 65 1002 158 1007
rect 385 1002 494 1007
rect 521 1002 750 1007
rect 817 1002 846 1007
rect 897 1002 902 1012
rect 2641 1007 2646 1032
rect 2665 1022 2806 1027
rect 2849 1022 2902 1027
rect 2665 1012 2742 1017
rect 2809 1012 2878 1017
rect 2897 1007 2902 1022
rect 961 1002 1006 1007
rect 1017 1002 1102 1007
rect 1681 1002 1702 1007
rect 1897 1002 2062 1007
rect 2641 1002 2686 1007
rect 2713 1002 2782 1007
rect 2873 1002 2902 1007
rect 961 997 966 1002
rect 1121 997 1342 1002
rect 161 992 286 997
rect 313 992 398 997
rect 537 992 638 997
rect 761 992 878 997
rect 889 992 966 997
rect 977 992 1126 997
rect 1337 992 1510 997
rect 1641 992 1670 997
rect 1689 992 1726 997
rect 1777 992 1950 997
rect 1969 992 2054 997
rect 2193 992 2238 997
rect 2569 992 2702 997
rect 2729 992 2910 997
rect 129 982 254 987
rect 265 982 438 987
rect 809 982 990 987
rect 1001 982 1326 987
rect 2025 982 2214 987
rect 2593 982 2670 987
rect 2793 982 2846 987
rect 2913 982 2950 987
rect 1369 977 1486 982
rect 177 972 206 977
rect 257 972 374 977
rect 905 972 1374 977
rect 1481 972 1510 977
rect 2617 972 2702 977
rect 2761 972 2926 977
rect 585 962 718 967
rect 737 962 982 967
rect 1097 962 1150 967
rect 1385 962 1518 967
rect 2017 962 2062 967
rect 2081 962 2126 967
rect 2625 962 2678 967
rect 2705 962 2742 967
rect 2801 962 2878 967
rect 585 957 590 962
rect 561 952 590 957
rect 713 957 718 962
rect 1169 957 1342 962
rect 713 952 750 957
rect 913 952 950 957
rect 1105 952 1174 957
rect 1337 952 1422 957
rect 1497 952 1582 957
rect 1881 952 2118 957
rect 2129 952 2150 957
rect 2497 952 2526 957
rect 2609 952 2854 957
rect 2881 952 2958 957
rect 2881 947 2886 952
rect 129 942 190 947
rect 385 942 526 947
rect 641 942 702 947
rect 721 942 790 947
rect 1057 942 1110 947
rect 1137 942 1326 947
rect 1497 942 1558 947
rect 1761 942 1822 947
rect 2073 942 2134 947
rect 2185 942 2246 947
rect 2473 942 2526 947
rect 2665 942 2742 947
rect 2753 942 2886 947
rect 2897 942 2934 947
rect 2961 942 2990 947
rect 385 937 390 942
rect 361 932 390 937
rect 521 937 526 942
rect 785 937 790 942
rect 521 932 662 937
rect 785 932 822 937
rect 889 932 926 937
rect 961 932 1022 937
rect 1289 932 1374 937
rect 1777 932 1894 937
rect 1041 927 1182 932
rect 81 922 246 927
rect 313 922 414 927
rect 513 922 614 927
rect 625 922 806 927
rect 825 922 918 927
rect 937 922 1046 927
rect 1177 922 1398 927
rect 1713 922 1766 927
rect 1785 922 1870 927
rect 177 912 230 917
rect 377 912 502 917
rect 697 912 758 917
rect 329 902 366 907
rect 569 902 654 907
rect 673 902 718 907
rect 569 897 574 902
rect 321 892 350 897
rect 345 887 350 892
rect 417 892 446 897
rect 481 892 574 897
rect 649 897 654 902
rect 801 897 806 922
rect 977 912 1094 917
rect 1121 912 1166 917
rect 1313 912 1526 917
rect 1601 912 1678 917
rect 1697 912 1750 917
rect 1777 912 1846 917
rect 1873 912 1902 917
rect 1601 907 1606 912
rect 913 902 958 907
rect 977 902 1030 907
rect 1297 902 1462 907
rect 1561 902 1606 907
rect 1673 907 1678 912
rect 2001 907 2006 937
rect 2489 932 2550 937
rect 2601 932 2718 937
rect 2049 922 2134 927
rect 2201 922 2342 927
rect 2417 922 2494 927
rect 2505 922 2614 927
rect 2721 922 2750 927
rect 2745 917 2750 922
rect 2849 922 2918 927
rect 2849 917 2854 922
rect 2393 912 2438 917
rect 2465 912 2494 917
rect 1673 902 1798 907
rect 2001 902 2158 907
rect 913 897 918 902
rect 2489 897 2494 912
rect 2689 912 2718 917
rect 2745 912 2854 917
rect 2913 917 2918 922
rect 2913 912 2966 917
rect 2689 897 2694 912
rect 2873 902 2974 907
rect 649 892 710 897
rect 801 892 918 897
rect 937 892 974 897
rect 1153 892 1246 897
rect 1385 892 1518 897
rect 1617 892 1782 897
rect 417 887 422 892
rect 1777 887 1782 892
rect 1913 892 2158 897
rect 2489 892 2694 897
rect 1913 887 1918 892
rect 345 882 422 887
rect 585 882 686 887
rect 1209 882 1238 887
rect 1233 877 1238 882
rect 1369 882 1398 887
rect 1665 882 1758 887
rect 1777 882 1918 887
rect 2225 882 2318 887
rect 1369 877 1374 882
rect 625 872 742 877
rect 1233 872 1374 877
rect 2761 872 2830 877
rect 1673 862 1726 867
rect 2345 862 2382 867
rect 2601 862 2662 867
rect 2889 862 2998 867
rect 473 852 710 857
rect 1441 852 1630 857
rect 2073 852 2174 857
rect 2361 852 2438 857
rect 2457 852 2518 857
rect 1441 847 1446 852
rect 1417 842 1446 847
rect 1625 847 1630 852
rect 1625 842 1750 847
rect 1929 842 1966 847
rect 2041 842 2166 847
rect 2193 842 2262 847
rect 2369 842 2726 847
rect 2193 837 2198 842
rect 361 832 414 837
rect 433 832 478 837
rect 601 832 686 837
rect 1081 832 1134 837
rect 1537 832 1614 837
rect 1969 832 2198 837
rect 2257 837 2262 842
rect 2721 837 2726 842
rect 2257 832 2334 837
rect 2385 832 2430 837
rect 2721 832 2750 837
rect 2897 832 2950 837
rect 2569 827 2638 832
rect 137 822 198 827
rect 393 822 550 827
rect 561 822 670 827
rect 777 822 838 827
rect 857 822 974 827
rect 1025 822 1118 827
rect 1393 822 1486 827
rect 1721 822 1758 827
rect 1993 822 2094 827
rect 2353 822 2382 827
rect 2521 822 2574 827
rect 2633 822 2870 827
rect 2921 822 2958 827
rect 545 817 550 822
rect 857 817 862 822
rect 185 812 214 817
rect 329 812 390 817
rect 417 812 526 817
rect 545 812 574 817
rect 585 812 614 817
rect 697 812 734 817
rect 793 812 862 817
rect 969 817 974 822
rect 969 812 1046 817
rect 209 807 214 812
rect 1041 807 1046 812
rect 1137 812 1166 817
rect 1209 812 1390 817
rect 1465 812 1702 817
rect 1881 812 2014 817
rect 2081 812 2126 817
rect 2145 812 2198 817
rect 2217 812 2246 817
rect 2385 812 2494 817
rect 2585 812 2622 817
rect 1137 807 1142 812
rect 1697 807 1702 812
rect 1793 807 1862 812
rect 2865 807 2870 822
rect 2889 812 2942 817
rect 193 802 214 807
rect 465 802 518 807
rect 585 802 686 807
rect 825 802 854 807
rect 1041 802 1142 807
rect 1233 802 1478 807
rect 1697 802 1798 807
rect 1857 802 2118 807
rect 2129 802 2174 807
rect 2345 802 2382 807
rect 2553 802 2614 807
rect 2689 802 2742 807
rect 2865 802 2942 807
rect 681 797 830 802
rect 185 792 246 797
rect 377 792 430 797
rect 561 792 630 797
rect 873 792 958 797
rect 1241 792 1350 797
rect 1497 792 1558 797
rect 1601 792 1630 797
rect 1657 792 1742 797
rect 1809 792 1870 797
rect 1985 792 2014 797
rect 2097 792 2150 797
rect 2225 792 2270 797
rect 2569 792 2678 797
rect 2857 792 2918 797
rect 129 782 182 787
rect 201 782 318 787
rect 353 782 406 787
rect 513 782 646 787
rect 729 782 1022 787
rect 1161 782 1278 787
rect 1369 782 1478 787
rect 1745 782 1854 787
rect 1985 782 2046 787
rect 2137 782 2182 787
rect 2201 782 2286 787
rect 2353 782 2398 787
rect 2665 782 2870 787
rect 2921 782 2990 787
rect 177 777 182 782
rect 1369 777 1374 782
rect 177 772 310 777
rect 361 772 438 777
rect 569 772 630 777
rect 641 772 798 777
rect 897 772 926 777
rect 217 762 358 767
rect 353 757 358 762
rect 449 762 502 767
rect 449 757 454 762
rect 297 752 334 757
rect 353 752 454 757
rect 497 757 502 762
rect 641 757 646 772
rect 921 767 926 772
rect 1025 772 1054 777
rect 1185 772 1374 777
rect 1473 777 1478 782
rect 1473 772 1558 777
rect 1737 772 1774 777
rect 1817 772 1878 777
rect 2097 772 2118 777
rect 2833 772 2974 777
rect 1025 767 1030 772
rect 721 762 894 767
rect 921 762 1030 767
rect 1049 762 1526 767
rect 1897 762 2054 767
rect 2441 762 2518 767
rect 2441 757 2446 762
rect 497 752 646 757
rect 721 752 886 757
rect 1169 752 1254 757
rect 1289 752 1422 757
rect 1417 747 1422 752
rect 1529 752 1718 757
rect 1753 752 1782 757
rect 1841 752 2046 757
rect 2409 752 2446 757
rect 2513 757 2518 762
rect 2513 752 2590 757
rect 2673 752 2742 757
rect 1529 747 1534 752
rect 1713 747 1718 752
rect 665 742 710 747
rect 745 742 806 747
rect 921 742 1022 747
rect 1145 742 1310 747
rect 1417 742 1534 747
rect 1553 742 1574 747
rect 1713 742 1758 747
rect 1105 732 1158 737
rect 1249 732 1286 737
rect 409 722 510 727
rect 529 722 598 727
rect 641 722 718 727
rect 889 722 926 727
rect 1009 722 1070 727
rect 1121 722 1238 727
rect 409 717 414 722
rect 169 712 342 717
rect 385 712 414 717
rect 505 717 510 722
rect 641 717 646 722
rect 505 712 550 717
rect 617 712 646 717
rect 713 717 718 722
rect 713 712 742 717
rect 761 712 870 717
rect 881 712 966 717
rect 1073 712 1134 717
rect 1305 712 1414 717
rect 1553 712 1558 742
rect 1569 732 1710 737
rect 1777 727 1782 752
rect 2737 747 2742 752
rect 1801 742 1910 747
rect 2025 742 2086 747
rect 2513 742 2582 747
rect 2681 742 2710 747
rect 2737 742 2766 747
rect 2785 742 2998 747
rect 1865 732 1982 737
rect 2161 732 2222 737
rect 2457 732 2494 737
rect 2049 727 2142 732
rect 1753 722 1782 727
rect 1841 722 2054 727
rect 2137 722 2414 727
rect 2705 722 2798 727
rect 2881 722 3006 727
rect 1593 712 1638 717
rect 1729 712 1758 717
rect 1305 707 1310 712
rect 289 702 342 707
rect 441 702 734 707
rect 1241 702 1310 707
rect 1409 707 1414 712
rect 1753 707 1758 712
rect 1849 712 1878 717
rect 1913 712 1942 717
rect 2065 712 2142 717
rect 2169 712 2286 717
rect 2537 712 2806 717
rect 2825 712 2902 717
rect 1849 707 1854 712
rect 2801 707 2806 712
rect 1409 702 1438 707
rect 1753 702 1854 707
rect 1881 702 1942 707
rect 2449 702 2534 707
rect 2801 702 2854 707
rect 417 692 534 697
rect 625 692 654 697
rect 649 687 654 692
rect 721 692 750 697
rect 1281 692 1614 697
rect 2809 692 2854 697
rect 721 687 726 692
rect 649 682 726 687
rect 1385 682 1422 687
rect 1889 682 2078 687
rect 2273 682 2334 687
rect 2513 672 2654 677
rect 505 662 614 667
rect 1897 662 1950 667
rect 505 657 510 662
rect 481 652 510 657
rect 609 657 614 662
rect 2513 657 2518 672
rect 609 652 638 657
rect 969 652 1110 657
rect 1313 652 1542 657
rect 1969 652 2062 657
rect 369 642 462 647
rect 369 637 374 642
rect 345 632 374 637
rect 457 637 462 642
rect 969 637 974 652
rect 457 632 622 637
rect 657 632 686 637
rect 945 632 974 637
rect 1105 637 1110 652
rect 1969 647 1974 652
rect 1945 642 1974 647
rect 2057 647 2062 652
rect 2105 652 2182 657
rect 2361 652 2390 657
rect 2489 652 2518 657
rect 2649 657 2654 672
rect 2649 652 2846 657
rect 2105 647 2110 652
rect 2057 642 2110 647
rect 2177 647 2182 652
rect 2177 642 2206 647
rect 2433 642 2462 647
rect 2481 642 2638 647
rect 1105 632 1238 637
rect 1313 632 1342 637
rect 1809 632 1886 637
rect 1937 632 2070 637
rect 2441 632 2510 637
rect 2689 632 2726 637
rect 2889 632 2942 637
rect 1313 627 1318 632
rect 1809 627 1814 632
rect 177 622 278 627
rect 297 622 494 627
rect 665 622 726 627
rect 769 622 878 627
rect 929 622 1038 627
rect 1057 622 1094 627
rect 1289 622 1318 627
rect 1353 622 1398 627
rect 1417 622 1510 627
rect 1529 622 1718 627
rect 1785 622 1814 627
rect 1881 627 1886 632
rect 1881 622 1910 627
rect 2121 622 2238 627
rect 2273 622 2398 627
rect 2417 622 2518 627
rect 2665 622 2726 627
rect 2865 622 2934 627
rect 1113 617 1270 622
rect 1417 617 1422 622
rect 225 612 294 617
rect 313 612 398 617
rect 425 612 462 617
rect 657 612 694 617
rect 857 612 1054 617
rect 1065 612 1118 617
rect 1265 612 1422 617
rect 1505 617 1510 622
rect 2273 617 2278 622
rect 1505 612 1558 617
rect 1801 612 1982 617
rect 2089 612 2126 617
rect 2249 612 2278 617
rect 2393 617 2398 622
rect 2393 612 2438 617
rect 2857 612 2902 617
rect 713 607 830 612
rect 1553 607 1558 612
rect 2121 607 2254 612
rect 185 602 326 607
rect 473 602 526 607
rect 625 602 718 607
rect 825 602 894 607
rect 913 602 974 607
rect 1105 602 1174 607
rect 1201 602 1518 607
rect 1553 602 1574 607
rect 2017 602 2102 607
rect 1201 597 1206 602
rect 2897 597 2902 612
rect 233 592 286 597
rect 401 592 502 597
rect 569 592 662 597
rect 729 592 814 597
rect 1025 592 1094 597
rect 1113 592 1206 597
rect 1217 592 1254 597
rect 1313 592 1342 597
rect 1457 592 1486 597
rect 1601 592 1646 597
rect 1761 592 1830 597
rect 1945 592 2006 597
rect 2105 592 2166 597
rect 2289 592 2374 597
rect 2417 592 2526 597
rect 2673 592 2774 597
rect 2897 592 2926 597
rect 161 582 246 587
rect 449 582 718 587
rect 929 582 1126 587
rect 1177 582 1438 587
rect 1489 582 1582 587
rect 1753 582 1806 587
rect 2065 582 2398 587
rect 2409 582 2430 587
rect 89 572 150 577
rect 145 567 150 572
rect 241 572 366 577
rect 417 572 470 577
rect 585 572 646 577
rect 985 572 1086 577
rect 1345 572 1526 577
rect 1593 572 1798 577
rect 2129 572 2190 577
rect 2273 572 2318 577
rect 241 567 246 572
rect 1105 567 1174 572
rect 1241 567 1326 572
rect 1521 567 1598 572
rect 145 562 246 567
rect 617 562 774 567
rect 849 562 950 567
rect 1049 562 1110 567
rect 1169 562 1246 567
rect 1321 562 1390 567
rect 1465 562 1502 567
rect 1961 562 2382 567
rect 2449 562 2566 567
rect 769 557 774 562
rect 265 552 302 557
rect 705 552 750 557
rect 769 552 1086 557
rect 1121 552 1158 557
rect 1257 552 1494 557
rect 1577 552 1606 557
rect 1617 552 1654 557
rect 1777 552 1926 557
rect 2145 552 2334 557
rect 2441 552 2494 557
rect 2873 552 2942 557
rect 1153 547 1262 552
rect 161 542 190 547
rect 305 542 446 547
rect 465 542 566 547
rect 697 542 758 547
rect 769 542 878 547
rect 945 542 982 547
rect 1073 542 1134 547
rect 1281 542 1414 547
rect 1425 542 1486 547
rect 1561 542 1590 547
rect 465 537 470 542
rect 137 532 158 537
rect 433 532 470 537
rect 561 537 566 542
rect 1585 537 1590 542
rect 1665 542 1734 547
rect 1937 542 1982 547
rect 2113 542 2174 547
rect 2425 542 2494 547
rect 2777 542 2934 547
rect 1665 537 1670 542
rect 561 532 662 537
rect 825 532 1030 537
rect 1041 532 1166 537
rect 1305 532 1334 537
rect 1393 532 1494 537
rect 1585 532 1670 537
rect 2105 532 2182 537
rect 2553 532 2606 537
rect 2649 532 2742 537
rect 401 522 534 527
rect 561 522 582 527
rect 833 522 886 527
rect 1017 522 1070 527
rect 1329 522 1358 527
rect 1425 522 1470 527
rect 1689 522 1742 527
rect 1905 522 2150 527
rect 2273 522 2358 527
rect 2465 522 2582 527
rect 2625 522 2710 527
rect 2945 522 2950 547
rect 1089 517 1206 522
rect 113 512 262 517
rect 417 512 638 517
rect 785 512 822 517
rect 1009 512 1030 517
rect 1041 512 1094 517
rect 1201 512 1302 517
rect 1329 512 1334 522
rect 1393 512 1438 517
rect 1553 512 1582 517
rect 1633 512 1678 517
rect 1857 512 1894 517
rect 2129 512 2246 517
rect 2617 512 2686 517
rect 2697 512 2790 517
rect 313 502 390 507
rect 489 502 582 507
rect 793 502 846 507
rect 1057 502 1190 507
rect 1441 502 1614 507
rect 2401 502 2430 507
rect 2905 502 2942 507
rect 569 492 726 497
rect 945 492 998 497
rect 993 487 998 492
rect 1177 492 1262 497
rect 1801 492 1878 497
rect 1897 492 1918 497
rect 2409 492 2446 497
rect 2561 492 2598 497
rect 1177 487 1182 492
rect 993 482 1182 487
rect 1201 482 1286 487
rect 2201 482 2254 487
rect 169 472 206 477
rect 2089 472 2222 477
rect 1953 462 2030 467
rect 1953 457 1958 462
rect 817 452 894 457
rect 913 452 1030 457
rect 1865 452 1958 457
rect 2025 457 2030 462
rect 2025 452 2054 457
rect 2385 452 2414 457
rect 817 447 822 452
rect 305 442 406 447
rect 577 442 702 447
rect 753 442 822 447
rect 889 447 894 452
rect 889 442 934 447
rect 1041 442 1070 447
rect 1529 442 1630 447
rect 1969 442 2110 447
rect 305 437 310 442
rect 281 432 310 437
rect 401 437 406 442
rect 929 437 1046 442
rect 401 432 486 437
rect 505 432 590 437
rect 713 432 766 437
rect 833 432 910 437
rect 1473 432 1526 437
rect 1569 432 1638 437
rect 1793 432 1846 437
rect 1993 432 2062 437
rect 2105 432 2286 437
rect 2457 432 2566 437
rect 1841 427 1846 432
rect 153 422 190 427
rect 273 422 342 427
rect 425 422 558 427
rect 625 422 742 427
rect 881 422 918 427
rect 913 417 918 422
rect 1001 422 1030 427
rect 1089 422 1134 427
rect 1537 422 1590 427
rect 1745 422 1790 427
rect 1841 422 1950 427
rect 2033 422 2086 427
rect 2273 422 2310 427
rect 2785 422 2822 427
rect 1001 417 1006 422
rect 1945 417 1950 422
rect 121 412 166 417
rect 321 412 486 417
rect 497 412 518 417
rect 569 412 614 417
rect 777 412 894 417
rect 913 412 1006 417
rect 1249 412 1270 417
rect 1425 412 1486 417
rect 1505 412 1534 417
rect 1593 412 1630 417
rect 1769 412 1822 417
rect 1945 412 2062 417
rect 2265 412 2294 417
rect 2713 412 2870 417
rect 1081 402 1182 407
rect 1617 402 1670 407
rect 1849 402 1934 407
rect 2065 402 2094 407
rect 2761 402 2846 407
rect 2913 402 2934 407
rect 1929 397 2070 402
rect 153 392 198 397
rect 209 392 238 397
rect 257 392 302 397
rect 377 392 534 397
rect 769 392 830 397
rect 1065 392 1134 397
rect 1257 392 1302 397
rect 1321 392 1454 397
rect 1737 392 1790 397
rect 1841 392 1886 397
rect 2105 392 2150 397
rect 2209 392 2294 397
rect 2313 392 2414 397
rect 2641 392 2734 397
rect 2913 392 2918 402
rect 2929 392 2966 397
rect 193 387 198 392
rect 1321 387 1326 392
rect 193 382 318 387
rect 385 382 510 387
rect 537 382 758 387
rect 785 382 942 387
rect 977 382 1326 387
rect 1449 387 1454 392
rect 2289 387 2294 392
rect 1449 382 1478 387
rect 1769 382 1990 387
rect 2289 382 2422 387
rect 2673 382 2742 387
rect 2881 382 2958 387
rect 129 372 214 377
rect 241 372 326 377
rect 737 372 798 377
rect 1105 372 1198 377
rect 1281 372 1814 377
rect 1913 372 2206 377
rect 2529 372 2926 377
rect 921 362 974 367
rect 1065 362 1094 367
rect 1817 362 1974 367
rect 2081 362 2126 367
rect 2249 362 2422 367
rect 2665 362 2726 367
rect 2897 362 2974 367
rect 1401 357 1502 362
rect 1969 357 2086 362
rect 281 352 414 357
rect 825 352 902 357
rect 937 352 982 357
rect 1025 352 1094 357
rect 1377 352 1406 357
rect 1497 352 1526 357
rect 1785 352 1910 357
rect 2705 352 2758 357
rect 825 347 830 352
rect 177 342 206 347
rect 329 342 390 347
rect 433 342 582 347
rect 601 342 646 347
rect 665 342 782 347
rect 801 342 830 347
rect 897 347 902 352
rect 897 342 950 347
rect 1033 342 1118 347
rect 1217 342 1278 347
rect 1409 342 1566 347
rect 1849 342 1934 347
rect 1953 342 2038 347
rect 2049 342 2078 347
rect 2193 342 2254 347
rect 2313 342 2438 347
rect 433 337 438 342
rect 161 332 294 337
rect 321 332 438 337
rect 577 337 582 342
rect 665 337 670 342
rect 577 332 670 337
rect 777 337 782 342
rect 777 332 1022 337
rect 1129 332 1214 337
rect 1233 332 1254 337
rect 1425 332 1454 337
rect 1609 332 1646 337
rect 1793 332 1862 337
rect 1921 332 2022 337
rect 2033 332 2062 337
rect 2153 332 2246 337
rect 2673 332 2814 337
rect 1017 327 1134 332
rect 145 322 206 327
rect 201 317 206 322
rect 305 322 334 327
rect 345 322 438 327
rect 537 322 574 327
rect 633 322 678 327
rect 697 322 782 327
rect 865 322 910 327
rect 1249 322 1254 332
rect 1281 322 1342 327
rect 1377 322 1422 327
rect 1449 322 1614 327
rect 1985 322 2014 327
rect 2433 322 2494 327
rect 305 317 310 322
rect 1281 317 1286 322
rect 81 312 182 317
rect 201 312 310 317
rect 449 312 502 317
rect 665 312 742 317
rect 809 312 1062 317
rect 1233 312 1286 317
rect 1345 312 1406 317
rect 1433 312 1470 317
rect 1553 312 1598 317
rect 1625 312 1678 317
rect 1905 312 1990 317
rect 1985 307 1990 312
rect 2073 312 2206 317
rect 2281 312 2358 317
rect 2513 312 2614 317
rect 2633 312 2918 317
rect 2073 307 2078 312
rect 2513 307 2518 312
rect 513 302 550 307
rect 593 302 710 307
rect 745 302 854 307
rect 889 302 926 307
rect 921 297 926 302
rect 1009 302 1038 307
rect 1353 302 1398 307
rect 1417 302 1598 307
rect 1857 302 1966 307
rect 1985 302 2078 307
rect 2441 302 2518 307
rect 2609 307 2614 312
rect 2609 302 2654 307
rect 2745 302 2774 307
rect 1009 297 1014 302
rect 2769 297 2774 302
rect 2841 302 2870 307
rect 2841 297 2846 302
rect 697 292 774 297
rect 833 292 902 297
rect 921 292 1014 297
rect 1337 292 1382 297
rect 1441 292 1470 297
rect 2497 292 2598 297
rect 2769 292 2846 297
rect 217 282 694 287
rect 713 282 862 287
rect 689 277 694 282
rect 689 272 1222 277
rect 1513 272 1654 277
rect 321 262 606 267
rect 673 262 718 267
rect 753 262 822 267
rect 2065 262 2230 267
rect 321 257 326 262
rect 297 252 326 257
rect 601 257 606 262
rect 2065 257 2070 262
rect 601 252 630 257
rect 841 252 926 257
rect 1425 252 1462 257
rect 1977 252 2070 257
rect 345 247 494 252
rect 729 247 846 252
rect 921 247 926 252
rect 1977 247 1982 252
rect 289 242 350 247
rect 489 242 678 247
rect 705 242 734 247
rect 921 242 950 247
rect 1473 242 1542 247
rect 1889 242 1982 247
rect 2225 247 2230 262
rect 2529 252 2630 257
rect 2529 247 2534 252
rect 2225 242 2254 247
rect 2505 242 2534 247
rect 2625 247 2630 252
rect 2625 242 2654 247
rect 201 232 350 237
rect 369 232 1134 237
rect 1377 232 1550 237
rect 369 227 374 232
rect 161 222 286 227
rect 329 222 374 227
rect 401 222 438 227
rect 505 222 566 227
rect 657 222 830 227
rect 865 222 910 227
rect 1105 222 1230 227
rect 1241 222 1358 227
rect 1441 222 1526 227
rect 209 212 318 217
rect 553 212 846 217
rect 889 212 918 217
rect 961 212 1054 217
rect 1393 212 1430 217
rect 1473 212 1574 217
rect 1585 212 1590 237
rect 2081 232 2174 237
rect 2233 232 2286 237
rect 2313 232 2342 237
rect 2497 232 2526 237
rect 2553 227 2678 232
rect 1881 222 1902 227
rect 1993 222 2110 227
rect 2161 222 2246 227
rect 2329 222 2382 227
rect 2529 222 2558 227
rect 2673 222 2702 227
rect 2761 222 2790 227
rect 2889 222 2926 227
rect 2241 217 2246 222
rect 1609 212 1638 217
rect 1833 212 1918 217
rect 1985 212 2054 217
rect 2241 212 2350 217
rect 2489 212 2518 217
rect 2545 212 2638 217
rect 401 207 534 212
rect 961 207 966 212
rect 177 202 254 207
rect 249 197 254 202
rect 329 202 406 207
rect 529 202 830 207
rect 937 202 966 207
rect 1049 207 1054 212
rect 1049 202 1182 207
rect 329 197 334 202
rect 825 197 942 202
rect 1473 197 1478 212
rect 1977 202 2038 207
rect 2681 202 2790 207
rect 1513 197 1622 202
rect 129 192 230 197
rect 249 192 334 197
rect 417 192 478 197
rect 537 192 694 197
rect 721 192 806 197
rect 977 192 1038 197
rect 1121 192 1214 197
rect 1225 192 1286 197
rect 1361 192 1478 197
rect 1489 192 1518 197
rect 1617 192 1646 197
rect 1913 192 1958 197
rect 2121 192 2182 197
rect 2321 192 2406 197
rect 2521 192 2590 197
rect 2705 192 2734 197
rect 2729 187 2734 192
rect 2801 192 2862 197
rect 2801 187 2806 192
rect 169 182 214 187
rect 449 182 1166 187
rect 1369 182 1606 187
rect 1945 182 1990 187
rect 2009 182 2086 187
rect 2361 182 2470 187
rect 2729 182 2806 187
rect 2889 182 2910 187
rect 449 177 454 182
rect 1225 177 1318 182
rect 201 172 270 177
rect 297 172 454 177
rect 473 172 614 177
rect 625 172 774 177
rect 1201 172 1230 177
rect 1313 172 1598 177
rect 1937 172 1982 177
rect 2345 172 2438 177
rect 273 162 310 167
rect 457 162 654 167
rect 833 162 910 167
rect 937 162 998 167
rect 1209 162 1366 167
rect 2273 162 2494 167
rect 2561 162 2766 167
rect 113 157 206 162
rect 329 157 438 162
rect 673 157 814 162
rect 89 152 118 157
rect 201 152 334 157
rect 433 152 678 157
rect 809 152 1262 157
rect 1329 152 1446 157
rect 2345 152 2382 157
rect 2529 152 2566 157
rect 2705 152 2838 157
rect 137 142 190 147
rect 257 142 614 147
rect 633 142 710 147
rect 769 142 886 147
rect 937 142 1030 147
rect 1153 142 1374 147
rect 1393 142 1462 147
rect 1785 142 1886 147
rect 2081 142 2198 147
rect 2329 142 2374 147
rect 2489 142 2558 147
rect 2673 142 2750 147
rect 2825 142 2942 147
rect 609 137 614 142
rect 425 132 486 137
rect 609 132 806 137
rect 1185 132 1270 137
rect 1449 132 1470 137
rect 2169 132 2318 137
rect 305 127 430 132
rect 2313 127 2318 132
rect 2393 132 2454 137
rect 2393 127 2398 132
rect 289 122 310 127
rect 449 122 742 127
rect 881 122 958 127
rect 1377 122 1486 127
rect 1561 122 1598 127
rect 2313 122 2398 127
rect 2457 122 2486 127
rect 2513 122 2894 127
rect 185 112 278 117
rect 385 112 470 117
rect 497 112 606 117
rect 641 112 702 117
rect 809 112 894 117
rect 985 112 1086 117
rect 1345 112 1406 117
rect 1449 112 1478 117
rect 2065 112 2158 117
rect 2153 107 2158 112
rect 2257 112 2286 117
rect 2473 112 2630 117
rect 2257 107 2262 112
rect 489 102 518 107
rect 513 87 518 102
rect 713 102 782 107
rect 1585 102 1622 107
rect 2153 102 2262 107
rect 2465 102 2494 107
rect 2505 102 2534 107
rect 713 87 718 102
rect 2529 97 2534 102
rect 2665 102 2694 107
rect 2921 102 2974 107
rect 2665 97 2670 102
rect 2529 92 2670 97
rect 513 82 718 87
<< gv2 >>
rect 3095 2863 3097 2865
rect 3095 2813 3097 2815
rect 3095 2733 3097 2735
rect 3095 2613 3097 2615
rect 3095 2533 3097 2535
rect 3095 2413 3097 2415
rect -4 2363 -2 2365
rect 3095 2363 3097 2365
rect -4 2293 -2 2295
rect 3095 2263 3097 2265
rect 3095 2183 3097 2185
rect 3095 2163 3097 2165
rect 3095 2143 3097 2145
rect -5 2013 -3 2015
rect 3095 2013 3097 2015
rect -5 1993 -3 1995
rect 3095 1933 3097 1935
rect -4 1923 -2 1925
rect 3095 1913 3097 1915
rect -4 1903 -2 1905
use Project_Top_VIA1  Project_Top_VIA1_0
timestamp 1681620392
transform 1 0 24 0 1 3017
box -10 -10 10 10
use M3_M2  M3_M2_0
timestamp 1681620392
transform 1 0 1852 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1681620392
transform 1 0 1884 0 1 3025
box -3 -3 3 3
use Project_Top_VIA1  Project_Top_VIA1_1
timestamp 1681620392
transform 1 0 3067 0 1 3017
box -10 -10 10 10
use Project_Top_VIA1  Project_Top_VIA1_2
timestamp 1681620392
transform 1 0 48 0 1 2993
box -10 -10 10 10
use M3_M2  M3_M2_2
timestamp 1681620392
transform 1 0 2228 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3
timestamp 1681620392
transform 1 0 2284 0 1 2995
box -3 -3 3 3
use Project_Top_VIA1  Project_Top_VIA1_3
timestamp 1681620392
transform 1 0 3043 0 1 2993
box -10 -10 10 10
use Project_Top_VIA0  Project_Top_VIA0_0
timestamp 1681620392
transform 1 0 48 0 1 2970
box -10 -3 10 3
use M3_M2  M3_M2_52
timestamp 1681620392
transform 1 0 84 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_2
timestamp 1681620392
transform 1 0 124 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_53
timestamp 1681620392
transform 1 0 124 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_56
timestamp 1681620392
transform 1 0 172 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_57
timestamp 1681620392
transform 1 0 204 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_58
timestamp 1681620392
transform 1 0 220 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_59
timestamp 1681620392
transform 1 0 236 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1681620392
transform 1 0 236 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_70
timestamp 1681620392
transform 1 0 244 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_60
timestamp 1681620392
transform 1 0 268 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_119
timestamp 1681620392
transform 1 0 252 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1681620392
transform 1 0 260 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_138
timestamp 1681620392
transform 1 0 244 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1681620392
transform 1 0 260 0 1 2905
box -2 -2 2 2
use M3_M2  M3_M2_86
timestamp 1681620392
transform 1 0 268 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1681620392
transform 1 0 324 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3
timestamp 1681620392
transform 1 0 316 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_54
timestamp 1681620392
transform 1 0 316 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_4
timestamp 1681620392
transform 1 0 340 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1681620392
transform 1 0 316 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1681620392
transform 1 0 332 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5
timestamp 1681620392
transform 1 0 364 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_61
timestamp 1681620392
transform 1 0 356 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_87
timestamp 1681620392
transform 1 0 332 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_88
timestamp 1681620392
transform 1 0 356 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_93
timestamp 1681620392
transform 1 0 340 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_62
timestamp 1681620392
transform 1 0 396 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_71
timestamp 1681620392
transform 1 0 404 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_43
timestamp 1681620392
transform 1 0 420 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_123
timestamp 1681620392
transform 1 0 412 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_94
timestamp 1681620392
transform 1 0 388 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_6
timestamp 1681620392
transform 1 0 460 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_44
timestamp 1681620392
transform 1 0 476 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_72
timestamp 1681620392
transform 1 0 476 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1681620392
transform 1 0 524 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1681620392
transform 1 0 540 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1681620392
transform 1 0 532 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_7
timestamp 1681620392
transform 1 0 532 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_8
timestamp 1681620392
transform 1 0 540 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_55
timestamp 1681620392
transform 1 0 516 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_63
timestamp 1681620392
transform 1 0 524 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_64
timestamp 1681620392
transform 1 0 540 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_124
timestamp 1681620392
transform 1 0 508 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_89
timestamp 1681620392
transform 1 0 508 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_9
timestamp 1681620392
transform 1 0 572 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_45
timestamp 1681620392
transform 1 0 580 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_10
timestamp 1681620392
transform 1 0 588 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_65
timestamp 1681620392
transform 1 0 564 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_56
timestamp 1681620392
transform 1 0 572 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_66
timestamp 1681620392
transform 1 0 580 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_67
timestamp 1681620392
transform 1 0 596 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_4
timestamp 1681620392
transform 1 0 604 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_18
timestamp 1681620392
transform 1 0 612 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_11
timestamp 1681620392
transform 1 0 604 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_12
timestamp 1681620392
transform 1 0 612 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_73
timestamp 1681620392
transform 1 0 564 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_74
timestamp 1681620392
transform 1 0 596 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_90
timestamp 1681620392
transform 1 0 564 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1681620392
transform 1 0 644 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_19
timestamp 1681620392
transform 1 0 636 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1681620392
transform 1 0 668 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_13
timestamp 1681620392
transform 1 0 628 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_14
timestamp 1681620392
transform 1 0 652 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_15
timestamp 1681620392
transform 1 0 668 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_68
timestamp 1681620392
transform 1 0 636 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_69
timestamp 1681620392
transform 1 0 644 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_57
timestamp 1681620392
transform 1 0 652 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_70
timestamp 1681620392
transform 1 0 660 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1681620392
transform 1 0 684 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_9
timestamp 1681620392
transform 1 0 692 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_16
timestamp 1681620392
transform 1 0 692 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_58
timestamp 1681620392
transform 1 0 700 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_125
timestamp 1681620392
transform 1 0 700 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_17
timestamp 1681620392
transform 1 0 716 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_5
timestamp 1681620392
transform 1 0 748 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_46
timestamp 1681620392
transform 1 0 764 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_72
timestamp 1681620392
transform 1 0 740 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_59
timestamp 1681620392
transform 1 0 748 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_73
timestamp 1681620392
transform 1 0 772 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_75
timestamp 1681620392
transform 1 0 740 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_60
timestamp 1681620392
transform 1 0 780 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_74
timestamp 1681620392
transform 1 0 788 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_61
timestamp 1681620392
transform 1 0 796 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_75
timestamp 1681620392
transform 1 0 804 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_126
timestamp 1681620392
transform 1 0 748 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_127
timestamp 1681620392
transform 1 0 756 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_140
timestamp 1681620392
transform 1 0 732 0 1 2905
box -2 -2 2 2
use M3_M2  M3_M2_76
timestamp 1681620392
transform 1 0 772 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_128
timestamp 1681620392
transform 1 0 780 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_77
timestamp 1681620392
transform 1 0 788 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_141
timestamp 1681620392
transform 1 0 764 0 1 2905
box -2 -2 2 2
use M3_M2  M3_M2_95
timestamp 1681620392
transform 1 0 732 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_96
timestamp 1681620392
transform 1 0 756 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_18
timestamp 1681620392
transform 1 0 820 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1681620392
transform 1 0 836 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_19
timestamp 1681620392
transform 1 0 860 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_21
timestamp 1681620392
transform 1 0 948 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_20
timestamp 1681620392
transform 1 0 972 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_77
timestamp 1681620392
transform 1 0 892 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_78
timestamp 1681620392
transform 1 0 948 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_78
timestamp 1681620392
transform 1 0 892 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_21
timestamp 1681620392
transform 1 0 988 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_79
timestamp 1681620392
transform 1 0 988 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_22
timestamp 1681620392
transform 1 0 1012 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_22
timestamp 1681620392
transform 1 0 1012 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_129
timestamp 1681620392
transform 1 0 1012 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_23
timestamp 1681620392
transform 1 0 1068 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_23
timestamp 1681620392
transform 1 0 1044 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_24
timestamp 1681620392
transform 1 0 1172 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_0
timestamp 1681620392
transform 1 0 1180 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_24
timestamp 1681620392
transform 1 0 1148 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_25
timestamp 1681620392
transform 1 0 1164 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_26
timestamp 1681620392
transform 1 0 1180 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_79
timestamp 1681620392
transform 1 0 1068 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_80
timestamp 1681620392
transform 1 0 1124 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_62
timestamp 1681620392
transform 1 0 1148 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_81
timestamp 1681620392
transform 1 0 1164 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_80
timestamp 1681620392
transform 1 0 1116 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_81
timestamp 1681620392
transform 1 0 1164 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_25
timestamp 1681620392
transform 1 0 1300 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_27
timestamp 1681620392
transform 1 0 1300 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_82
timestamp 1681620392
transform 1 0 1204 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1681620392
transform 1 0 1212 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_84
timestamp 1681620392
transform 1 0 1220 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_85
timestamp 1681620392
transform 1 0 1268 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_63
timestamp 1681620392
transform 1 0 1300 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_26
timestamp 1681620392
transform 1 0 1316 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_28
timestamp 1681620392
transform 1 0 1332 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_64
timestamp 1681620392
transform 1 0 1332 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_27
timestamp 1681620392
transform 1 0 1476 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_29
timestamp 1681620392
transform 1 0 1428 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1681620392
transform 1 0 1356 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1681620392
transform 1 0 1412 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_88
timestamp 1681620392
transform 1 0 1476 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_89
timestamp 1681620392
transform 1 0 1508 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_28
timestamp 1681620392
transform 1 0 1540 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_30
timestamp 1681620392
transform 1 0 1540 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_130
timestamp 1681620392
transform 1 0 1540 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_31
timestamp 1681620392
transform 1 0 1580 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_90
timestamp 1681620392
transform 1 0 1564 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1681620392
transform 1 0 1572 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1
timestamp 1681620392
transform 1 0 1612 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_32
timestamp 1681620392
transform 1 0 1604 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_33
timestamp 1681620392
transform 1 0 1644 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1681620392
transform 1 0 1644 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_29
timestamp 1681620392
transform 1 0 1684 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_30
timestamp 1681620392
transform 1 0 1724 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_34
timestamp 1681620392
transform 1 0 1684 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_35
timestamp 1681620392
transform 1 0 1772 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_92
timestamp 1681620392
transform 1 0 1660 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1681620392
transform 1 0 1668 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_65
timestamp 1681620392
transform 1 0 1676 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_94
timestamp 1681620392
transform 1 0 1692 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_66
timestamp 1681620392
transform 1 0 1708 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_95
timestamp 1681620392
transform 1 0 1724 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1681620392
transform 1 0 1684 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_82
timestamp 1681620392
transform 1 0 1740 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_83
timestamp 1681620392
transform 1 0 1772 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_97
timestamp 1681620392
transform 1 0 1692 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_98
timestamp 1681620392
transform 1 0 1716 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_14
timestamp 1681620392
transform 1 0 1804 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_36
timestamp 1681620392
transform 1 0 1804 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_96
timestamp 1681620392
transform 1 0 1828 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_97
timestamp 1681620392
transform 1 0 1884 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_6
timestamp 1681620392
transform 1 0 1916 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_15
timestamp 1681620392
transform 1 0 1908 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_10
timestamp 1681620392
transform 1 0 1924 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_37
timestamp 1681620392
transform 1 0 1924 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_67
timestamp 1681620392
transform 1 0 1924 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_38
timestamp 1681620392
transform 1 0 2012 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_98
timestamp 1681620392
transform 1 0 1972 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1681620392
transform 1 0 2004 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_7
timestamp 1681620392
transform 1 0 2068 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_31
timestamp 1681620392
transform 1 0 2052 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_32
timestamp 1681620392
transform 1 0 2092 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_39
timestamp 1681620392
transform 1 0 2028 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_47
timestamp 1681620392
transform 1 0 2036 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_40
timestamp 1681620392
transform 1 0 2052 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_41
timestamp 1681620392
transform 1 0 2068 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_42
timestamp 1681620392
transform 1 0 2156 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_100
timestamp 1681620392
transform 1 0 2028 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_101
timestamp 1681620392
transform 1 0 2092 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_133
timestamp 1681620392
transform 1 0 2052 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_91
timestamp 1681620392
transform 1 0 2052 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_48
timestamp 1681620392
transform 1 0 2164 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_33
timestamp 1681620392
transform 1 0 2212 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_43
timestamp 1681620392
transform 1 0 2172 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_102
timestamp 1681620392
transform 1 0 2164 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_49
timestamp 1681620392
transform 1 0 2196 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_103
timestamp 1681620392
transform 1 0 2188 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1681620392
transform 1 0 2172 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_84
timestamp 1681620392
transform 1 0 2180 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_92
timestamp 1681620392
transform 1 0 2164 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1681620392
transform 1 0 2268 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_35
timestamp 1681620392
transform 1 0 2316 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_44
timestamp 1681620392
transform 1 0 2212 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_45
timestamp 1681620392
transform 1 0 2228 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_46
timestamp 1681620392
transform 1 0 2316 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_85
timestamp 1681620392
transform 1 0 2204 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_135
timestamp 1681620392
transform 1 0 2212 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1681620392
transform 1 0 2268 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_36
timestamp 1681620392
transform 1 0 2348 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_47
timestamp 1681620392
transform 1 0 2348 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1681620392
transform 1 0 2380 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_106
timestamp 1681620392
transform 1 0 2428 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_37
timestamp 1681620392
transform 1 0 2524 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_48
timestamp 1681620392
transform 1 0 2524 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1681620392
transform 1 0 2444 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_108
timestamp 1681620392
transform 1 0 2500 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_38
timestamp 1681620392
transform 1 0 2556 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_49
timestamp 1681620392
transform 1 0 2556 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1681620392
transform 1 0 2580 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_110
timestamp 1681620392
transform 1 0 2636 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_39
timestamp 1681620392
transform 1 0 2668 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_50
timestamp 1681620392
transform 1 0 2668 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_51
timestamp 1681620392
transform 1 0 2756 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_111
timestamp 1681620392
transform 1 0 2700 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_40
timestamp 1681620392
transform 1 0 2860 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_50
timestamp 1681620392
transform 1 0 2780 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_51
timestamp 1681620392
transform 1 0 2820 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_52
timestamp 1681620392
transform 1 0 2860 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_112
timestamp 1681620392
transform 1 0 2764 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_113
timestamp 1681620392
transform 1 0 2780 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_114
timestamp 1681620392
transform 1 0 2836 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_68
timestamp 1681620392
transform 1 0 2860 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_136
timestamp 1681620392
transform 1 0 2772 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_53
timestamp 1681620392
transform 1 0 2884 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1681620392
transform 1 0 2876 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_69
timestamp 1681620392
transform 1 0 2884 0 1 2925
box -3 -3 3 3
use Project_Top_VIA0  Project_Top_VIA0_1
timestamp 1681620392
transform 1 0 3043 0 1 2970
box -10 -3 10 3
use M3_M2  M3_M2_16
timestamp 1681620392
transform 1 0 2932 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_41
timestamp 1681620392
transform 1 0 2916 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_42
timestamp 1681620392
transform 1 0 2956 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_54
timestamp 1681620392
transform 1 0 2916 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_55
timestamp 1681620392
transform 1 0 2932 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1681620392
transform 1 0 2956 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_117
timestamp 1681620392
transform 1 0 3012 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_137
timestamp 1681620392
transform 1 0 2916 0 1 2915
box -2 -2 2 2
use Project_Top_VIA0  Project_Top_VIA0_2
timestamp 1681620392
transform 1 0 24 0 1 2870
box -10 -3 10 3
use FILL  FILL_0
timestamp 1681620392
transform 1 0 72 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1
timestamp 1681620392
transform 1 0 80 0 -1 2970
box -8 -3 16 105
use FILL  FILL_2
timestamp 1681620392
transform 1 0 88 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3
timestamp 1681620392
transform 1 0 96 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4
timestamp 1681620392
transform 1 0 104 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_0
timestamp 1681620392
transform 1 0 112 0 -1 2970
box -8 -3 104 105
use FILL  FILL_5
timestamp 1681620392
transform 1 0 208 0 -1 2970
box -8 -3 16 105
use FILL  FILL_6
timestamp 1681620392
transform 1 0 216 0 -1 2970
box -8 -3 16 105
use NAND3X1  NAND3X1_0
timestamp 1681620392
transform 1 0 224 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_1
timestamp 1681620392
transform 1 0 256 0 -1 2970
box -8 -3 40 105
use FILL  FILL_7
timestamp 1681620392
transform 1 0 288 0 -1 2970
box -8 -3 16 105
use FILL  FILL_8
timestamp 1681620392
transform 1 0 296 0 -1 2970
box -8 -3 16 105
use FILL  FILL_9
timestamp 1681620392
transform 1 0 304 0 -1 2970
box -8 -3 16 105
use NAND2X1  NAND2X1_0
timestamp 1681620392
transform 1 0 312 0 -1 2970
box -8 -3 32 105
use OAI21X1  OAI21X1_0
timestamp 1681620392
transform -1 0 368 0 -1 2970
box -8 -3 34 105
use INVX2  INVX2_0
timestamp 1681620392
transform 1 0 368 0 -1 2970
box -9 -3 26 105
use OAI21X1  OAI21X1_1
timestamp 1681620392
transform 1 0 384 0 -1 2970
box -8 -3 34 105
use FILL  FILL_10
timestamp 1681620392
transform 1 0 416 0 -1 2970
box -8 -3 16 105
use FILL  FILL_11
timestamp 1681620392
transform 1 0 424 0 -1 2970
box -8 -3 16 105
use FILL  FILL_12
timestamp 1681620392
transform 1 0 432 0 -1 2970
box -8 -3 16 105
use FILL  FILL_13
timestamp 1681620392
transform 1 0 440 0 -1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_0
timestamp 1681620392
transform 1 0 448 0 -1 2970
box -8 -3 32 105
use FILL  FILL_14
timestamp 1681620392
transform 1 0 472 0 -1 2970
box -8 -3 16 105
use FILL  FILL_15
timestamp 1681620392
transform 1 0 480 0 -1 2970
box -8 -3 16 105
use FILL  FILL_16
timestamp 1681620392
transform 1 0 488 0 -1 2970
box -8 -3 16 105
use FILL  FILL_17
timestamp 1681620392
transform 1 0 496 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_2
timestamp 1681620392
transform -1 0 536 0 -1 2970
box -8 -3 34 105
use INVX2  INVX2_1
timestamp 1681620392
transform 1 0 536 0 -1 2970
box -9 -3 26 105
use OAI22X1  OAI22X1_0
timestamp 1681620392
transform 1 0 552 0 -1 2970
box -8 -3 46 105
use INVX2  INVX2_2
timestamp 1681620392
transform -1 0 608 0 -1 2970
box -9 -3 26 105
use FILL  FILL_18
timestamp 1681620392
transform 1 0 608 0 -1 2970
box -8 -3 16 105
use FILL  FILL_19
timestamp 1681620392
transform 1 0 616 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_3
timestamp 1681620392
transform 1 0 624 0 -1 2970
box -9 -3 26 105
use AOI22X1  AOI22X1_0
timestamp 1681620392
transform 1 0 640 0 -1 2970
box -8 -3 46 105
use INVX2  INVX2_4
timestamp 1681620392
transform -1 0 696 0 -1 2970
box -9 -3 26 105
use FILL  FILL_20
timestamp 1681620392
transform 1 0 696 0 -1 2970
box -8 -3 16 105
use FILL  FILL_21
timestamp 1681620392
transform 1 0 704 0 -1 2970
box -8 -3 16 105
use FILL  FILL_22
timestamp 1681620392
transform 1 0 712 0 -1 2970
box -8 -3 16 105
use NAND3X1  NAND3X1_2
timestamp 1681620392
transform -1 0 752 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_3
timestamp 1681620392
transform -1 0 784 0 -1 2970
box -8 -3 40 105
use INVX2  INVX2_5
timestamp 1681620392
transform -1 0 800 0 -1 2970
box -9 -3 26 105
use FILL  FILL_23
timestamp 1681620392
transform 1 0 800 0 -1 2970
box -8 -3 16 105
use FILL  FILL_24
timestamp 1681620392
transform 1 0 808 0 -1 2970
box -8 -3 16 105
use FILL  FILL_25
timestamp 1681620392
transform 1 0 816 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_6
timestamp 1681620392
transform -1 0 840 0 -1 2970
box -9 -3 26 105
use FILL  FILL_26
timestamp 1681620392
transform 1 0 840 0 -1 2970
box -8 -3 16 105
use FILL  FILL_27
timestamp 1681620392
transform 1 0 848 0 -1 2970
box -8 -3 16 105
use FILL  FILL_28
timestamp 1681620392
transform 1 0 856 0 -1 2970
box -8 -3 16 105
use FILL  FILL_29
timestamp 1681620392
transform 1 0 864 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_7
timestamp 1681620392
transform -1 0 888 0 -1 2970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_1
timestamp 1681620392
transform -1 0 984 0 -1 2970
box -8 -3 104 105
use FILL  FILL_30
timestamp 1681620392
transform 1 0 984 0 -1 2970
box -8 -3 16 105
use NAND2X1  NAND2X1_1
timestamp 1681620392
transform 1 0 992 0 -1 2970
box -8 -3 32 105
use OAI21X1  OAI21X1_3
timestamp 1681620392
transform -1 0 1048 0 -1 2970
box -8 -3 34 105
use INVX2  INVX2_8
timestamp 1681620392
transform -1 0 1064 0 -1 2970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_2
timestamp 1681620392
transform -1 0 1160 0 -1 2970
box -8 -3 104 105
use INVX2  INVX2_9
timestamp 1681620392
transform 1 0 1160 0 -1 2970
box -9 -3 26 105
use NOR2X1  NOR2X1_1
timestamp 1681620392
transform 1 0 1176 0 -1 2970
box -8 -3 32 105
use INVX2  INVX2_10
timestamp 1681620392
transform 1 0 1200 0 -1 2970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_3
timestamp 1681620392
transform -1 0 1312 0 -1 2970
box -8 -3 104 105
use FILL  FILL_31
timestamp 1681620392
transform 1 0 1312 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_4
timestamp 1681620392
transform 1 0 1320 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_5
timestamp 1681620392
transform 1 0 1416 0 -1 2970
box -8 -3 104 105
use FILL  FILL_32
timestamp 1681620392
transform 1 0 1512 0 -1 2970
box -8 -3 16 105
use NAND2X1  NAND2X1_2
timestamp 1681620392
transform 1 0 1520 0 -1 2970
box -8 -3 32 105
use OAI21X1  OAI21X1_4
timestamp 1681620392
transform -1 0 1576 0 -1 2970
box -8 -3 34 105
use FILL  FILL_33
timestamp 1681620392
transform 1 0 1576 0 -1 2970
box -8 -3 16 105
use OR2X1  OR2X1_0
timestamp 1681620392
transform -1 0 1616 0 -1 2970
box -8 -3 40 105
use FILL  FILL_34
timestamp 1681620392
transform 1 0 1616 0 -1 2970
box -8 -3 16 105
use NAND2X1  NAND2X1_3
timestamp 1681620392
transform 1 0 1624 0 -1 2970
box -8 -3 32 105
use FILL  FILL_35
timestamp 1681620392
transform 1 0 1648 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_5
timestamp 1681620392
transform 1 0 1656 0 -1 2970
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_6
timestamp 1681620392
transform -1 0 1784 0 -1 2970
box -8 -3 104 105
use FILL  FILL_36
timestamp 1681620392
transform 1 0 1784 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1681620392
transform 1 0 1792 0 -1 2970
box -8 -3 104 105
use FILL  FILL_37
timestamp 1681620392
transform 1 0 1888 0 -1 2970
box -8 -3 16 105
use FILL  FILL_38
timestamp 1681620392
transform 1 0 1896 0 -1 2970
box -8 -3 16 105
use FILL  FILL_39
timestamp 1681620392
transform 1 0 1904 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_8
timestamp 1681620392
transform 1 0 1912 0 -1 2970
box -8 -3 104 105
use FILL  FILL_40
timestamp 1681620392
transform 1 0 2008 0 -1 2970
box -8 -3 16 105
use FILL  FILL_41
timestamp 1681620392
transform 1 0 2016 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_6
timestamp 1681620392
transform 1 0 2024 0 -1 2970
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_9
timestamp 1681620392
transform 1 0 2056 0 -1 2970
box -8 -3 104 105
use NAND2X1  NAND2X1_4
timestamp 1681620392
transform 1 0 2152 0 -1 2970
box -8 -3 32 105
use OAI21X1  OAI21X1_7
timestamp 1681620392
transform 1 0 2176 0 -1 2970
box -8 -3 34 105
use NAND2X1  NAND2X1_5
timestamp 1681620392
transform -1 0 2232 0 -1 2970
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_10
timestamp 1681620392
transform -1 0 2328 0 -1 2970
box -8 -3 104 105
use FILL  FILL_42
timestamp 1681620392
transform 1 0 2328 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1681620392
transform 1 0 2336 0 -1 2970
box -8 -3 104 105
use FILL  FILL_43
timestamp 1681620392
transform 1 0 2432 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_12
timestamp 1681620392
transform -1 0 2536 0 -1 2970
box -8 -3 104 105
use FILL  FILL_44
timestamp 1681620392
transform 1 0 2536 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_13
timestamp 1681620392
transform 1 0 2544 0 -1 2970
box -8 -3 104 105
use FILL  FILL_45
timestamp 1681620392
transform 1 0 2640 0 -1 2970
box -8 -3 16 105
use FILL  FILL_46
timestamp 1681620392
transform 1 0 2648 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_14
timestamp 1681620392
transform 1 0 2656 0 -1 2970
box -8 -3 104 105
use NAND2X1  NAND2X1_6
timestamp 1681620392
transform 1 0 2752 0 -1 2970
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_15
timestamp 1681620392
transform -1 0 2872 0 -1 2970
box -8 -3 104 105
use FILL  FILL_47
timestamp 1681620392
transform 1 0 2872 0 -1 2970
box -8 -3 16 105
use FILL  FILL_48
timestamp 1681620392
transform 1 0 2880 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_8
timestamp 1681620392
transform 1 0 2888 0 -1 2970
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1681620392
transform 1 0 2920 0 -1 2970
box -8 -3 104 105
use Project_Top_VIA0  Project_Top_VIA0_3
timestamp 1681620392
transform 1 0 3067 0 1 2870
box -10 -3 10 3
use M2_M1  M2_M1_142
timestamp 1681620392
transform 1 0 116 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_143
timestamp 1681620392
transform 1 0 140 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_149
timestamp 1681620392
transform 1 0 124 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_144
timestamp 1681620392
transform 1 0 132 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_107
timestamp 1681620392
transform 1 0 172 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_144
timestamp 1681620392
transform 1 0 172 0 1 2835
box -2 -2 2 2
use M3_M2  M3_M2_117
timestamp 1681620392
transform 1 0 180 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_150
timestamp 1681620392
transform 1 0 148 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_151
timestamp 1681620392
transform 1 0 156 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_145
timestamp 1681620392
transform 1 0 164 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_152
timestamp 1681620392
transform 1 0 180 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_194
timestamp 1681620392
transform 1 0 132 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_203
timestamp 1681620392
transform 1 0 124 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_172
timestamp 1681620392
transform 1 0 148 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_195
timestamp 1681620392
transform 1 0 164 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_108
timestamp 1681620392
transform 1 0 212 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_196
timestamp 1681620392
transform 1 0 196 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_173
timestamp 1681620392
transform 1 0 204 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_276
timestamp 1681620392
transform 1 0 188 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_204
timestamp 1681620392
transform 1 0 196 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_277
timestamp 1681620392
transform 1 0 204 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_197
timestamp 1681620392
transform 1 0 236 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_278
timestamp 1681620392
transform 1 0 244 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_227
timestamp 1681620392
transform 1 0 236 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_145
timestamp 1681620392
transform 1 0 260 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_146
timestamp 1681620392
transform 1 0 276 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_153
timestamp 1681620392
transform 1 0 260 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1681620392
transform 1 0 268 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_198
timestamp 1681620392
transform 1 0 252 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_199
timestamp 1681620392
transform 1 0 268 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_205
timestamp 1681620392
transform 1 0 268 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_118
timestamp 1681620392
transform 1 0 292 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_206
timestamp 1681620392
transform 1 0 300 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_362
timestamp 1681620392
transform 1 0 292 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_155
timestamp 1681620392
transform 1 0 316 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_207
timestamp 1681620392
transform 1 0 316 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_279
timestamp 1681620392
transform 1 0 324 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_363
timestamp 1681620392
transform 1 0 324 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_156
timestamp 1681620392
transform 1 0 348 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1681620392
transform 1 0 340 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_208
timestamp 1681620392
transform 1 0 340 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_146
timestamp 1681620392
transform 1 0 372 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_201
timestamp 1681620392
transform 1 0 372 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_280
timestamp 1681620392
transform 1 0 364 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_228
timestamp 1681620392
transform 1 0 364 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_119
timestamp 1681620392
transform 1 0 404 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_147
timestamp 1681620392
transform 1 0 396 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_148
timestamp 1681620392
transform 1 0 412 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_202
timestamp 1681620392
transform 1 0 396 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_203
timestamp 1681620392
transform 1 0 412 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_281
timestamp 1681620392
transform 1 0 388 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1681620392
transform 1 0 404 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_283
timestamp 1681620392
transform 1 0 412 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_149
timestamp 1681620392
transform 1 0 452 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_204
timestamp 1681620392
transform 1 0 428 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_205
timestamp 1681620392
transform 1 0 436 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_364
timestamp 1681620392
transform 1 0 436 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_206
timestamp 1681620392
transform 1 0 460 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_209
timestamp 1681620392
transform 1 0 460 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_157
timestamp 1681620392
transform 1 0 476 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1681620392
transform 1 0 484 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_150
timestamp 1681620392
transform 1 0 508 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_174
timestamp 1681620392
transform 1 0 500 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_284
timestamp 1681620392
transform 1 0 500 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_285
timestamp 1681620392
transform 1 0 508 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_158
timestamp 1681620392
transform 1 0 524 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_175
timestamp 1681620392
transform 1 0 524 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_208
timestamp 1681620392
transform 1 0 532 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_210
timestamp 1681620392
transform 1 0 524 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_159
timestamp 1681620392
transform 1 0 540 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_151
timestamp 1681620392
transform 1 0 556 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_160
timestamp 1681620392
transform 1 0 572 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_176
timestamp 1681620392
transform 1 0 540 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_209
timestamp 1681620392
transform 1 0 556 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_210
timestamp 1681620392
transform 1 0 564 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1681620392
transform 1 0 540 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_287
timestamp 1681620392
transform 1 0 564 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_229
timestamp 1681620392
transform 1 0 532 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_177
timestamp 1681620392
transform 1 0 580 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_211
timestamp 1681620392
transform 1 0 588 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_178
timestamp 1681620392
transform 1 0 596 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_211
timestamp 1681620392
transform 1 0 588 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_253
timestamp 1681620392
transform 1 0 564 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_179
timestamp 1681620392
transform 1 0 620 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_288
timestamp 1681620392
transform 1 0 612 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_230
timestamp 1681620392
transform 1 0 604 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_212
timestamp 1681620392
transform 1 0 620 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_152
timestamp 1681620392
transform 1 0 636 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_212
timestamp 1681620392
transform 1 0 636 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_213
timestamp 1681620392
transform 1 0 644 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_289
timestamp 1681620392
transform 1 0 628 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_290
timestamp 1681620392
transform 1 0 636 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_365
timestamp 1681620392
transform 1 0 620 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_231
timestamp 1681620392
transform 1 0 636 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_254
timestamp 1681620392
transform 1 0 644 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_120
timestamp 1681620392
transform 1 0 668 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_153
timestamp 1681620392
transform 1 0 692 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_214
timestamp 1681620392
transform 1 0 676 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1681620392
transform 1 0 692 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_291
timestamp 1681620392
transform 1 0 684 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_161
timestamp 1681620392
transform 1 0 732 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1681620392
transform 1 0 716 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_154
timestamp 1681620392
transform 1 0 748 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_217
timestamp 1681620392
transform 1 0 740 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_292
timestamp 1681620392
transform 1 0 732 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_255
timestamp 1681620392
transform 1 0 740 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_121
timestamp 1681620392
transform 1 0 764 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_109
timestamp 1681620392
transform 1 0 780 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_110
timestamp 1681620392
transform 1 0 820 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_147
timestamp 1681620392
transform 1 0 796 0 1 2835
box -2 -2 2 2
use M3_M2  M3_M2_122
timestamp 1681620392
transform 1 0 820 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_148
timestamp 1681620392
transform 1 0 828 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_162
timestamp 1681620392
transform 1 0 772 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_293
timestamp 1681620392
transform 1 0 764 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_155
timestamp 1681620392
transform 1 0 788 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_163
timestamp 1681620392
transform 1 0 796 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_164
timestamp 1681620392
transform 1 0 820 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_218
timestamp 1681620392
transform 1 0 788 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_180
timestamp 1681620392
transform 1 0 796 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_219
timestamp 1681620392
transform 1 0 804 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_156
timestamp 1681620392
transform 1 0 836 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_165
timestamp 1681620392
transform 1 0 844 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_220
timestamp 1681620392
transform 1 0 836 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_294
timestamp 1681620392
transform 1 0 812 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_181
timestamp 1681620392
transform 1 0 844 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_157
timestamp 1681620392
transform 1 0 900 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_221
timestamp 1681620392
transform 1 0 900 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_222
timestamp 1681620392
transform 1 0 956 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_295
timestamp 1681620392
transform 1 0 980 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_232
timestamp 1681620392
transform 1 0 956 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_158
timestamp 1681620392
transform 1 0 996 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_123
timestamp 1681620392
transform 1 0 1012 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_166
timestamp 1681620392
transform 1 0 1020 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_167
timestamp 1681620392
transform 1 0 1028 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_182
timestamp 1681620392
transform 1 0 1004 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_223
timestamp 1681620392
transform 1 0 1012 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1681620392
transform 1 0 996 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_183
timestamp 1681620392
transform 1 0 1028 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_124
timestamp 1681620392
transform 1 0 1060 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_168
timestamp 1681620392
transform 1 0 1060 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_224
timestamp 1681620392
transform 1 0 1044 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_297
timestamp 1681620392
transform 1 0 1020 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_184
timestamp 1681620392
transform 1 0 1060 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_111
timestamp 1681620392
transform 1 0 1092 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_185
timestamp 1681620392
transform 1 0 1084 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_298
timestamp 1681620392
transform 1 0 1052 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1681620392
transform 1 0 1060 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_213
timestamp 1681620392
transform 1 0 1068 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_300
timestamp 1681620392
transform 1 0 1084 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_233
timestamp 1681620392
transform 1 0 1060 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_256
timestamp 1681620392
transform 1 0 1044 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_125
timestamp 1681620392
transform 1 0 1108 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_225
timestamp 1681620392
transform 1 0 1108 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_226
timestamp 1681620392
transform 1 0 1116 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_301
timestamp 1681620392
transform 1 0 1108 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_112
timestamp 1681620392
transform 1 0 1148 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_169
timestamp 1681620392
transform 1 0 1140 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_227
timestamp 1681620392
transform 1 0 1140 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1681620392
transform 1 0 1164 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1681620392
transform 1 0 1180 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1681620392
transform 1 0 1132 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_214
timestamp 1681620392
transform 1 0 1140 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_303
timestamp 1681620392
transform 1 0 1156 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_304
timestamp 1681620392
transform 1 0 1172 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_305
timestamp 1681620392
transform 1 0 1180 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_234
timestamp 1681620392
transform 1 0 1156 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_235
timestamp 1681620392
transform 1 0 1180 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_113
timestamp 1681620392
transform 1 0 1212 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_126
timestamp 1681620392
transform 1 0 1196 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_127
timestamp 1681620392
transform 1 0 1220 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_170
timestamp 1681620392
transform 1 0 1196 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_159
timestamp 1681620392
transform 1 0 1204 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_186
timestamp 1681620392
transform 1 0 1196 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_160
timestamp 1681620392
transform 1 0 1236 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_230
timestamp 1681620392
transform 1 0 1212 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_231
timestamp 1681620392
transform 1 0 1220 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_187
timestamp 1681620392
transform 1 0 1228 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_232
timestamp 1681620392
transform 1 0 1236 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_188
timestamp 1681620392
transform 1 0 1244 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_233
timestamp 1681620392
transform 1 0 1252 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_306
timestamp 1681620392
transform 1 0 1228 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_171
timestamp 1681620392
transform 1 0 1260 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_307
timestamp 1681620392
transform 1 0 1268 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_114
timestamp 1681620392
transform 1 0 1276 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_115
timestamp 1681620392
transform 1 0 1292 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_234
timestamp 1681620392
transform 1 0 1292 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1681620392
transform 1 0 1292 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1681620392
transform 1 0 1300 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_215
timestamp 1681620392
transform 1 0 1308 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_310
timestamp 1681620392
transform 1 0 1324 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_236
timestamp 1681620392
transform 1 0 1292 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_257
timestamp 1681620392
transform 1 0 1300 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_237
timestamp 1681620392
transform 1 0 1324 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_116
timestamp 1681620392
transform 1 0 1340 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_172
timestamp 1681620392
transform 1 0 1332 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_128
timestamp 1681620392
transform 1 0 1364 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_235
timestamp 1681620392
transform 1 0 1364 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_236
timestamp 1681620392
transform 1 0 1372 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1681620392
transform 1 0 1348 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_366
timestamp 1681620392
transform 1 0 1340 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_258
timestamp 1681620392
transform 1 0 1332 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_216
timestamp 1681620392
transform 1 0 1372 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_259
timestamp 1681620392
transform 1 0 1372 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_99
timestamp 1681620392
transform 1 0 1460 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_100
timestamp 1681620392
transform 1 0 1500 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_129
timestamp 1681620392
transform 1 0 1412 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_130
timestamp 1681620392
transform 1 0 1508 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_237
timestamp 1681620392
transform 1 0 1468 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_238
timestamp 1681620392
transform 1 0 1500 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_312
timestamp 1681620392
transform 1 0 1420 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_217
timestamp 1681620392
transform 1 0 1468 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_218
timestamp 1681620392
transform 1 0 1492 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_131
timestamp 1681620392
transform 1 0 1524 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_173
timestamp 1681620392
transform 1 0 1524 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1681620392
transform 1 0 1524 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_132
timestamp 1681620392
transform 1 0 1540 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_313
timestamp 1681620392
transform 1 0 1540 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1681620392
transform 1 0 1532 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_368
timestamp 1681620392
transform 1 0 1548 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_174
timestamp 1681620392
transform 1 0 1588 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_189
timestamp 1681620392
transform 1 0 1564 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_240
timestamp 1681620392
transform 1 0 1572 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_314
timestamp 1681620392
transform 1 0 1564 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_161
timestamp 1681620392
transform 1 0 1620 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1681620392
transform 1 0 1636 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_175
timestamp 1681620392
transform 1 0 1644 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_241
timestamp 1681620392
transform 1 0 1612 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_315
timestamp 1681620392
transform 1 0 1596 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_238
timestamp 1681620392
transform 1 0 1580 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_219
timestamp 1681620392
transform 1 0 1612 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_316
timestamp 1681620392
transform 1 0 1620 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1681620392
transform 1 0 1628 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_190
timestamp 1681620392
transform 1 0 1652 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_176
timestamp 1681620392
transform 1 0 1684 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_242
timestamp 1681620392
transform 1 0 1660 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_243
timestamp 1681620392
transform 1 0 1668 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_244
timestamp 1681620392
transform 1 0 1684 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1681620392
transform 1 0 1644 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_220
timestamp 1681620392
transform 1 0 1668 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_319
timestamp 1681620392
transform 1 0 1692 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_221
timestamp 1681620392
transform 1 0 1700 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_245
timestamp 1681620392
transform 1 0 1708 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1681620392
transform 1 0 1708 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_321
timestamp 1681620392
transform 1 0 1716 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_260
timestamp 1681620392
transform 1 0 1708 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_246
timestamp 1681620392
transform 1 0 1724 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_247
timestamp 1681620392
transform 1 0 1764 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_248
timestamp 1681620392
transform 1 0 1820 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_322
timestamp 1681620392
transform 1 0 1740 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_222
timestamp 1681620392
transform 1 0 1764 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_323
timestamp 1681620392
transform 1 0 1828 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_261
timestamp 1681620392
transform 1 0 1756 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_262
timestamp 1681620392
transform 1 0 1820 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_177
timestamp 1681620392
transform 1 0 1836 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_249
timestamp 1681620392
transform 1 0 1852 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_250
timestamp 1681620392
transform 1 0 1860 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_324
timestamp 1681620392
transform 1 0 1860 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_325
timestamp 1681620392
transform 1 0 1868 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_239
timestamp 1681620392
transform 1 0 1860 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_133
timestamp 1681620392
transform 1 0 1884 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_178
timestamp 1681620392
transform 1 0 1884 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_251
timestamp 1681620392
transform 1 0 1900 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_326
timestamp 1681620392
transform 1 0 1884 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_240
timestamp 1681620392
transform 1 0 1884 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_134
timestamp 1681620392
transform 1 0 1940 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_179
timestamp 1681620392
transform 1 0 1940 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_327
timestamp 1681620392
transform 1 0 1916 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_328
timestamp 1681620392
transform 1 0 1924 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_329
timestamp 1681620392
transform 1 0 1940 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_241
timestamp 1681620392
transform 1 0 1940 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_252
timestamp 1681620392
transform 1 0 1972 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_330
timestamp 1681620392
transform 1 0 1988 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1681620392
transform 1 0 2004 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_135
timestamp 1681620392
transform 1 0 2020 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_180
timestamp 1681620392
transform 1 0 2020 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_103
timestamp 1681620392
transform 1 0 2068 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_136
timestamp 1681620392
transform 1 0 2060 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_253
timestamp 1681620392
transform 1 0 2036 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_332
timestamp 1681620392
transform 1 0 2028 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_242
timestamp 1681620392
transform 1 0 2012 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_243
timestamp 1681620392
transform 1 0 2028 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_181
timestamp 1681620392
transform 1 0 2060 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_333
timestamp 1681620392
transform 1 0 2060 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_244
timestamp 1681620392
transform 1 0 2060 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_104
timestamp 1681620392
transform 1 0 2172 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_137
timestamp 1681620392
transform 1 0 2180 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_163
timestamp 1681620392
transform 1 0 2172 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_254
timestamp 1681620392
transform 1 0 2092 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_255
timestamp 1681620392
transform 1 0 2124 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1681620392
transform 1 0 2172 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_245
timestamp 1681620392
transform 1 0 2124 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_191
timestamp 1681620392
transform 1 0 2196 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_335
timestamp 1681620392
transform 1 0 2196 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_138
timestamp 1681620392
transform 1 0 2236 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_256
timestamp 1681620392
transform 1 0 2212 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_182
timestamp 1681620392
transform 1 0 2236 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_164
timestamp 1681620392
transform 1 0 2316 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_165
timestamp 1681620392
transform 1 0 2340 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_257
timestamp 1681620392
transform 1 0 2252 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_258
timestamp 1681620392
transform 1 0 2292 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_336
timestamp 1681620392
transform 1 0 2236 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_246
timestamp 1681620392
transform 1 0 2236 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_192
timestamp 1681620392
transform 1 0 2356 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1681620392
transform 1 0 2388 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_259
timestamp 1681620392
transform 1 0 2364 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1681620392
transform 1 0 2340 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_338
timestamp 1681620392
transform 1 0 2356 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_247
timestamp 1681620392
transform 1 0 2292 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_183
timestamp 1681620392
transform 1 0 2388 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_339
timestamp 1681620392
transform 1 0 2380 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_260
timestamp 1681620392
transform 1 0 2412 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_223
timestamp 1681620392
transform 1 0 2412 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_340
timestamp 1681620392
transform 1 0 2420 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_140
timestamp 1681620392
transform 1 0 2452 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_341
timestamp 1681620392
transform 1 0 2436 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_342
timestamp 1681620392
transform 1 0 2444 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1681620392
transform 1 0 2460 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_193
timestamp 1681620392
transform 1 0 2460 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_185
timestamp 1681620392
transform 1 0 2492 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_261
timestamp 1681620392
transform 1 0 2468 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_262
timestamp 1681620392
transform 1 0 2476 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_343
timestamp 1681620392
transform 1 0 2460 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_224
timestamp 1681620392
transform 1 0 2476 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_248
timestamp 1681620392
transform 1 0 2460 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_344
timestamp 1681620392
transform 1 0 2500 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_186
timestamp 1681620392
transform 1 0 2524 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_194
timestamp 1681620392
transform 1 0 2524 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_263
timestamp 1681620392
transform 1 0 2540 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_345
timestamp 1681620392
transform 1 0 2524 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_195
timestamp 1681620392
transform 1 0 2548 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_346
timestamp 1681620392
transform 1 0 2556 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_249
timestamp 1681620392
transform 1 0 2556 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_166
timestamp 1681620392
transform 1 0 2580 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_187
timestamp 1681620392
transform 1 0 2588 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_141
timestamp 1681620392
transform 1 0 2612 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_188
timestamp 1681620392
transform 1 0 2612 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_264
timestamp 1681620392
transform 1 0 2572 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_265
timestamp 1681620392
transform 1 0 2588 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_196
timestamp 1681620392
transform 1 0 2596 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_266
timestamp 1681620392
transform 1 0 2604 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_225
timestamp 1681620392
transform 1 0 2580 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_347
timestamp 1681620392
transform 1 0 2588 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_189
timestamp 1681620392
transform 1 0 2636 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_197
timestamp 1681620392
transform 1 0 2636 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_167
timestamp 1681620392
transform 1 0 2660 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_267
timestamp 1681620392
transform 1 0 2652 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_348
timestamp 1681620392
transform 1 0 2604 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_349
timestamp 1681620392
transform 1 0 2628 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_350
timestamp 1681620392
transform 1 0 2636 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_250
timestamp 1681620392
transform 1 0 2636 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_105
timestamp 1681620392
transform 1 0 2692 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_106
timestamp 1681620392
transform 1 0 2764 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_142
timestamp 1681620392
transform 1 0 2772 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_190
timestamp 1681620392
transform 1 0 2692 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_268
timestamp 1681620392
transform 1 0 2676 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_351
timestamp 1681620392
transform 1 0 2660 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_352
timestamp 1681620392
transform 1 0 2668 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_263
timestamp 1681620392
transform 1 0 2628 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_264
timestamp 1681620392
transform 1 0 2652 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_198
timestamp 1681620392
transform 1 0 2692 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_199
timestamp 1681620392
transform 1 0 2708 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_269
timestamp 1681620392
transform 1 0 2732 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_353
timestamp 1681620392
transform 1 0 2692 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_354
timestamp 1681620392
transform 1 0 2708 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_226
timestamp 1681620392
transform 1 0 2732 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_143
timestamp 1681620392
transform 1 0 2828 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_168
timestamp 1681620392
transform 1 0 2804 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_191
timestamp 1681620392
transform 1 0 2828 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_270
timestamp 1681620392
transform 1 0 2804 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_200
timestamp 1681620392
transform 1 0 2828 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_271
timestamp 1681620392
transform 1 0 2852 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_355
timestamp 1681620392
transform 1 0 2796 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_356
timestamp 1681620392
transform 1 0 2812 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1681620392
transform 1 0 2836 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_169
timestamp 1681620392
transform 1 0 2868 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_192
timestamp 1681620392
transform 1 0 2876 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_201
timestamp 1681620392
transform 1 0 2876 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_101
timestamp 1681620392
transform 1 0 2908 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_170
timestamp 1681620392
transform 1 0 2892 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_193
timestamp 1681620392
transform 1 0 2900 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_272
timestamp 1681620392
transform 1 0 2884 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_358
timestamp 1681620392
transform 1 0 2868 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_251
timestamp 1681620392
transform 1 0 2860 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_202
timestamp 1681620392
transform 1 0 2900 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_359
timestamp 1681620392
transform 1 0 2892 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_102
timestamp 1681620392
transform 1 0 3012 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_171
timestamp 1681620392
transform 1 0 3012 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_273
timestamp 1681620392
transform 1 0 2916 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_274
timestamp 1681620392
transform 1 0 2956 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_275
timestamp 1681620392
transform 1 0 3012 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1681620392
transform 1 0 2916 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_361
timestamp 1681620392
transform 1 0 2932 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_252
timestamp 1681620392
transform 1 0 2956 0 1 2795
box -3 -3 3 3
use Project_Top_VIA0  Project_Top_VIA0_4
timestamp 1681620392
transform 1 0 48 0 1 2770
box -10 -3 10 3
use FILL  FILL_49
timestamp 1681620392
transform 1 0 72 0 1 2770
box -8 -3 16 105
use FILL  FILL_51
timestamp 1681620392
transform 1 0 80 0 1 2770
box -8 -3 16 105
use FILL  FILL_53
timestamp 1681620392
transform 1 0 88 0 1 2770
box -8 -3 16 105
use FILL  FILL_55
timestamp 1681620392
transform 1 0 96 0 1 2770
box -8 -3 16 105
use FILL  FILL_57
timestamp 1681620392
transform 1 0 104 0 1 2770
box -8 -3 16 105
use FILL  FILL_59
timestamp 1681620392
transform 1 0 112 0 1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_4
timestamp 1681620392
transform 1 0 120 0 1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_5
timestamp 1681620392
transform 1 0 152 0 1 2770
box -8 -3 40 105
use INVX2  INVX2_11
timestamp 1681620392
transform 1 0 184 0 1 2770
box -9 -3 26 105
use FILL  FILL_60
timestamp 1681620392
transform 1 0 200 0 1 2770
box -8 -3 16 105
use FILL  FILL_61
timestamp 1681620392
transform 1 0 208 0 1 2770
box -8 -3 16 105
use FILL  FILL_62
timestamp 1681620392
transform 1 0 216 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_12
timestamp 1681620392
transform 1 0 224 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_13
timestamp 1681620392
transform 1 0 240 0 1 2770
box -9 -3 26 105
use NAND3X1  NAND3X1_6
timestamp 1681620392
transform 1 0 256 0 1 2770
box -8 -3 40 105
use FILL  FILL_63
timestamp 1681620392
transform 1 0 288 0 1 2770
box -8 -3 16 105
use FILL  FILL_64
timestamp 1681620392
transform 1 0 296 0 1 2770
box -8 -3 16 105
use FILL  FILL_65
timestamp 1681620392
transform 1 0 304 0 1 2770
box -8 -3 16 105
use FILL  FILL_66
timestamp 1681620392
transform 1 0 312 0 1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_2
timestamp 1681620392
transform 1 0 320 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_7
timestamp 1681620392
transform -1 0 368 0 1 2770
box -8 -3 32 105
use FILL  FILL_67
timestamp 1681620392
transform 1 0 368 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_1
timestamp 1681620392
transform 1 0 376 0 1 2770
box -8 -3 46 105
use INVX2  INVX2_14
timestamp 1681620392
transform 1 0 416 0 1 2770
box -9 -3 26 105
use AOI21X1  AOI21X1_0
timestamp 1681620392
transform -1 0 464 0 1 2770
box -7 -3 39 105
use FILL  FILL_68
timestamp 1681620392
transform 1 0 464 0 1 2770
box -8 -3 16 105
use NAND2X1  NAND2X1_8
timestamp 1681620392
transform -1 0 496 0 1 2770
box -8 -3 32 105
use FILL  FILL_69
timestamp 1681620392
transform 1 0 496 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_15
timestamp 1681620392
transform 1 0 504 0 1 2770
box -9 -3 26 105
use FILL  FILL_70
timestamp 1681620392
transform 1 0 520 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_265
timestamp 1681620392
transform 1 0 540 0 1 2775
box -3 -3 3 3
use FILL  FILL_71
timestamp 1681620392
transform 1 0 528 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_266
timestamp 1681620392
transform 1 0 572 0 1 2775
box -3 -3 3 3
use OAI21X1  OAI21X1_9
timestamp 1681620392
transform -1 0 568 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_10
timestamp 1681620392
transform -1 0 600 0 1 2770
box -8 -3 34 105
use FILL  FILL_72
timestamp 1681620392
transform 1 0 600 0 1 2770
box -8 -3 16 105
use FILL  FILL_73
timestamp 1681620392
transform 1 0 608 0 1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_3
timestamp 1681620392
transform 1 0 616 0 1 2770
box -8 -3 32 105
use FILL  FILL_74
timestamp 1681620392
transform 1 0 640 0 1 2770
box -8 -3 16 105
use FILL  FILL_75
timestamp 1681620392
transform 1 0 648 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_2
timestamp 1681620392
transform 1 0 656 0 1 2770
box -8 -3 46 105
use FILL  FILL_76
timestamp 1681620392
transform 1 0 696 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_11
timestamp 1681620392
transform 1 0 704 0 1 2770
box -8 -3 34 105
use INVX2  INVX2_16
timestamp 1681620392
transform -1 0 752 0 1 2770
box -9 -3 26 105
use FILL  FILL_77
timestamp 1681620392
transform 1 0 752 0 1 2770
box -8 -3 16 105
use FILL  FILL_78
timestamp 1681620392
transform 1 0 760 0 1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_7
timestamp 1681620392
transform -1 0 800 0 1 2770
box -8 -3 40 105
use INVX2  INVX2_17
timestamp 1681620392
transform -1 0 816 0 1 2770
box -9 -3 26 105
use M3_M2  M3_M2_267
timestamp 1681620392
transform 1 0 828 0 1 2775
box -3 -3 3 3
use NAND3X1  NAND3X1_8
timestamp 1681620392
transform -1 0 848 0 1 2770
box -8 -3 40 105
use FILL  FILL_79
timestamp 1681620392
transform 1 0 848 0 1 2770
box -8 -3 16 105
use FILL  FILL_80
timestamp 1681620392
transform 1 0 856 0 1 2770
box -8 -3 16 105
use FILL  FILL_81
timestamp 1681620392
transform 1 0 864 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_268
timestamp 1681620392
transform 1 0 892 0 1 2775
box -3 -3 3 3
use INVX2  INVX2_18
timestamp 1681620392
transform -1 0 888 0 1 2770
box -9 -3 26 105
use FILL  FILL_82
timestamp 1681620392
transform 1 0 888 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_269
timestamp 1681620392
transform 1 0 988 0 1 2775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_17
timestamp 1681620392
transform -1 0 992 0 1 2770
box -8 -3 104 105
use FILL  FILL_83
timestamp 1681620392
transform 1 0 992 0 1 2770
box -8 -3 16 105
use NAND2X1  NAND2X1_9
timestamp 1681620392
transform 1 0 1000 0 1 2770
box -8 -3 32 105
use OAI21X1  OAI21X1_12
timestamp 1681620392
transform -1 0 1056 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_13
timestamp 1681620392
transform -1 0 1088 0 1 2770
box -8 -3 34 105
use FILL  FILL_84
timestamp 1681620392
transform 1 0 1088 0 1 2770
box -8 -3 16 105
use FILL  FILL_85
timestamp 1681620392
transform 1 0 1096 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_14
timestamp 1681620392
transform 1 0 1104 0 1 2770
box -8 -3 34 105
use FILL  FILL_86
timestamp 1681620392
transform 1 0 1136 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_270
timestamp 1681620392
transform 1 0 1172 0 1 2775
box -3 -3 3 3
use AOI22X1  AOI22X1_3
timestamp 1681620392
transform -1 0 1184 0 1 2770
box -8 -3 46 105
use FILL  FILL_87
timestamp 1681620392
transform 1 0 1184 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_15
timestamp 1681620392
transform -1 0 1224 0 1 2770
box -8 -3 34 105
use M3_M2  M3_M2_271
timestamp 1681620392
transform 1 0 1260 0 1 2775
box -3 -3 3 3
use OAI21X1  OAI21X1_16
timestamp 1681620392
transform 1 0 1224 0 1 2770
box -8 -3 34 105
use FILL  FILL_88
timestamp 1681620392
transform 1 0 1256 0 1 2770
box -8 -3 16 105
use FILL  FILL_89
timestamp 1681620392
transform 1 0 1264 0 1 2770
box -8 -3 16 105
use FILL  FILL_100
timestamp 1681620392
transform 1 0 1272 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_24
timestamp 1681620392
transform -1 0 1296 0 1 2770
box -9 -3 26 105
use OAI21X1  OAI21X1_22
timestamp 1681620392
transform 1 0 1296 0 1 2770
box -8 -3 34 105
use M3_M2  M3_M2_272
timestamp 1681620392
transform 1 0 1340 0 1 2775
box -3 -3 3 3
use FILL  FILL_101
timestamp 1681620392
transform 1 0 1328 0 1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_8
timestamp 1681620392
transform 1 0 1336 0 1 2770
box -8 -3 32 105
use INVX2  INVX2_25
timestamp 1681620392
transform 1 0 1360 0 1 2770
box -9 -3 26 105
use FILL  FILL_102
timestamp 1681620392
transform 1 0 1376 0 1 2770
box -8 -3 16 105
use FILL  FILL_103
timestamp 1681620392
transform 1 0 1384 0 1 2770
box -8 -3 16 105
use FILL  FILL_107
timestamp 1681620392
transform 1 0 1392 0 1 2770
box -8 -3 16 105
use FILL  FILL_108
timestamp 1681620392
transform 1 0 1400 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_22
timestamp 1681620392
transform 1 0 1408 0 1 2770
box -8 -3 104 105
use NAND2X1  NAND2X1_13
timestamp 1681620392
transform 1 0 1504 0 1 2770
box -8 -3 32 105
use FILL  FILL_109
timestamp 1681620392
transform 1 0 1528 0 1 2770
box -8 -3 16 105
use FILL  FILL_112
timestamp 1681620392
transform 1 0 1536 0 1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_9
timestamp 1681620392
transform 1 0 1544 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_14
timestamp 1681620392
transform 1 0 1568 0 1 2770
box -8 -3 32 105
use OAI21X1  OAI21X1_25
timestamp 1681620392
transform -1 0 1624 0 1 2770
box -8 -3 34 105
use M3_M2  M3_M2_273
timestamp 1681620392
transform 1 0 1644 0 1 2775
box -3 -3 3 3
use NAND2X1  NAND2X1_15
timestamp 1681620392
transform 1 0 1624 0 1 2770
box -8 -3 32 105
use FILL  FILL_113
timestamp 1681620392
transform 1 0 1648 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_26
timestamp 1681620392
transform 1 0 1656 0 1 2770
box -8 -3 34 105
use FILL  FILL_114
timestamp 1681620392
transform 1 0 1688 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_274
timestamp 1681620392
transform 1 0 1716 0 1 2775
box -3 -3 3 3
use INVX2  INVX2_26
timestamp 1681620392
transform -1 0 1712 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_27
timestamp 1681620392
transform 1 0 1712 0 1 2770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_24
timestamp 1681620392
transform 1 0 1728 0 1 2770
box -8 -3 104 105
use FILL  FILL_115
timestamp 1681620392
transform 1 0 1824 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_27
timestamp 1681620392
transform -1 0 1864 0 1 2770
box -8 -3 34 105
use NAND2X1  NAND2X1_16
timestamp 1681620392
transform 1 0 1864 0 1 2770
box -8 -3 32 105
use OAI21X1  OAI21X1_28
timestamp 1681620392
transform 1 0 1888 0 1 2770
box -8 -3 34 105
use NAND2X1  NAND2X1_17
timestamp 1681620392
transform 1 0 1920 0 1 2770
box -8 -3 32 105
use FILL  FILL_116
timestamp 1681620392
transform 1 0 1944 0 1 2770
box -8 -3 16 105
use FILL  FILL_117
timestamp 1681620392
transform 1 0 1952 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_29
timestamp 1681620392
transform 1 0 1960 0 1 2770
box -8 -3 34 105
use FILL  FILL_118
timestamp 1681620392
transform 1 0 1992 0 1 2770
box -8 -3 16 105
use NAND2X1  NAND2X1_18
timestamp 1681620392
transform 1 0 2000 0 1 2770
box -8 -3 32 105
use OAI21X1  OAI21X1_30
timestamp 1681620392
transform 1 0 2024 0 1 2770
box -8 -3 34 105
use NAND2X1  NAND2X1_19
timestamp 1681620392
transform -1 0 2080 0 1 2770
box -8 -3 32 105
use FILL  FILL_119
timestamp 1681620392
transform 1 0 2080 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_25
timestamp 1681620392
transform -1 0 2184 0 1 2770
box -8 -3 104 105
use FILL  FILL_120
timestamp 1681620392
transform 1 0 2184 0 1 2770
box -8 -3 16 105
use FILL  FILL_121
timestamp 1681620392
transform 1 0 2192 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_31
timestamp 1681620392
transform 1 0 2200 0 1 2770
box -8 -3 34 105
use NAND2X1  NAND2X1_20
timestamp 1681620392
transform -1 0 2256 0 1 2770
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_26
timestamp 1681620392
transform -1 0 2352 0 1 2770
box -8 -3 104 105
use OAI21X1  OAI21X1_32
timestamp 1681620392
transform 1 0 2352 0 1 2770
box -8 -3 34 105
use NAND2X1  NAND2X1_21
timestamp 1681620392
transform -1 0 2408 0 1 2770
box -8 -3 32 105
use FILL  FILL_122
timestamp 1681620392
transform 1 0 2408 0 1 2770
box -8 -3 16 105
use FILL  FILL_123
timestamp 1681620392
transform 1 0 2416 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_28
timestamp 1681620392
transform -1 0 2440 0 1 2770
box -9 -3 26 105
use NAND2X1  NAND2X1_22
timestamp 1681620392
transform 1 0 2440 0 1 2770
box -8 -3 32 105
use OAI21X1  OAI21X1_33
timestamp 1681620392
transform 1 0 2464 0 1 2770
box -8 -3 34 105
use FILL  FILL_124
timestamp 1681620392
transform 1 0 2496 0 1 2770
box -8 -3 16 105
use FILL  FILL_125
timestamp 1681620392
transform 1 0 2504 0 1 2770
box -8 -3 16 105
use FILL  FILL_126
timestamp 1681620392
transform 1 0 2512 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_34
timestamp 1681620392
transform -1 0 2552 0 1 2770
box -8 -3 34 105
use FILL  FILL_127
timestamp 1681620392
transform 1 0 2552 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_35
timestamp 1681620392
transform 1 0 2560 0 1 2770
box -8 -3 34 105
use INVX2  INVX2_29
timestamp 1681620392
transform -1 0 2608 0 1 2770
box -9 -3 26 105
use NAND2X1  NAND2X1_23
timestamp 1681620392
transform -1 0 2632 0 1 2770
box -8 -3 32 105
use M3_M2  M3_M2_275
timestamp 1681620392
transform 1 0 2652 0 1 2775
box -3 -3 3 3
use OAI21X1  OAI21X1_36
timestamp 1681620392
transform -1 0 2664 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_37
timestamp 1681620392
transform 1 0 2664 0 1 2770
box -8 -3 34 105
use M3_M2  M3_M2_276
timestamp 1681620392
transform 1 0 2708 0 1 2775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_27
timestamp 1681620392
transform 1 0 2696 0 1 2770
box -8 -3 104 105
use INVX2  INVX2_30
timestamp 1681620392
transform 1 0 2792 0 1 2770
box -9 -3 26 105
use NAND2X1  NAND2X1_24
timestamp 1681620392
transform 1 0 2808 0 1 2770
box -8 -3 32 105
use OAI21X1  OAI21X1_38
timestamp 1681620392
transform -1 0 2864 0 1 2770
box -8 -3 34 105
use FILL  FILL_128
timestamp 1681620392
transform 1 0 2864 0 1 2770
box -8 -3 16 105
use NAND2X1  NAND2X1_25
timestamp 1681620392
transform -1 0 2896 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_26
timestamp 1681620392
transform -1 0 2920 0 1 2770
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_28
timestamp 1681620392
transform 1 0 2920 0 1 2770
box -8 -3 104 105
use Project_Top_VIA0  Project_Top_VIA0_5
timestamp 1681620392
transform 1 0 3043 0 1 2770
box -10 -3 10 3
use M3_M2  M3_M2_399
timestamp 1681620392
transform 1 0 84 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_286
timestamp 1681620392
transform 1 0 116 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_376
timestamp 1681620392
transform 1 0 148 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_442
timestamp 1681620392
transform 1 0 124 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_443
timestamp 1681620392
transform 1 0 148 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_523
timestamp 1681620392
transform 1 0 116 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_369
timestamp 1681620392
transform 1 0 172 0 1 2745
box -2 -2 2 2
use M3_M2  M3_M2_333
timestamp 1681620392
transform 1 0 172 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_444
timestamp 1681620392
transform 1 0 172 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_524
timestamp 1681620392
transform 1 0 140 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_550
timestamp 1681620392
transform 1 0 132 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_382
timestamp 1681620392
transform 1 0 156 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_433
timestamp 1681620392
transform 1 0 140 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_287
timestamp 1681620392
transform 1 0 188 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_288
timestamp 1681620392
transform 1 0 244 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_289
timestamp 1681620392
transform 1 0 292 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_370
timestamp 1681620392
transform 1 0 188 0 1 2745
box -2 -2 2 2
use M3_M2  M3_M2_305
timestamp 1681620392
transform 1 0 276 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_377
timestamp 1681620392
transform 1 0 188 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_334
timestamp 1681620392
transform 1 0 196 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_335
timestamp 1681620392
transform 1 0 244 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_378
timestamp 1681620392
transform 1 0 276 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_360
timestamp 1681620392
transform 1 0 188 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_445
timestamp 1681620392
transform 1 0 196 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_446
timestamp 1681620392
transform 1 0 244 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_383
timestamp 1681620392
transform 1 0 180 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_371
timestamp 1681620392
transform 1 0 324 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_447
timestamp 1681620392
transform 1 0 300 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_361
timestamp 1681620392
transform 1 0 308 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_525
timestamp 1681620392
transform 1 0 292 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_400
timestamp 1681620392
transform 1 0 276 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_401
timestamp 1681620392
transform 1 0 292 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_290
timestamp 1681620392
transform 1 0 348 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_291
timestamp 1681620392
transform 1 0 364 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_292
timestamp 1681620392
transform 1 0 388 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_293
timestamp 1681620392
transform 1 0 404 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_306
timestamp 1681620392
transform 1 0 380 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_379
timestamp 1681620392
transform 1 0 332 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_380
timestamp 1681620392
transform 1 0 340 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_336
timestamp 1681620392
transform 1 0 348 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_381
timestamp 1681620392
transform 1 0 364 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_337
timestamp 1681620392
transform 1 0 372 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_382
timestamp 1681620392
transform 1 0 380 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_338
timestamp 1681620392
transform 1 0 388 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_307
timestamp 1681620392
transform 1 0 420 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_372
timestamp 1681620392
transform 1 0 428 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_383
timestamp 1681620392
transform 1 0 404 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_384
timestamp 1681620392
transform 1 0 412 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_362
timestamp 1681620392
transform 1 0 332 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_448
timestamp 1681620392
transform 1 0 340 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_449
timestamp 1681620392
transform 1 0 364 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_450
timestamp 1681620392
transform 1 0 372 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_451
timestamp 1681620392
transform 1 0 388 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_452
timestamp 1681620392
transform 1 0 404 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_526
timestamp 1681620392
transform 1 0 316 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_551
timestamp 1681620392
transform 1 0 308 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_418
timestamp 1681620392
transform 1 0 212 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_419
timestamp 1681620392
transform 1 0 284 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_420
timestamp 1681620392
transform 1 0 316 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_402
timestamp 1681620392
transform 1 0 340 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_403
timestamp 1681620392
transform 1 0 364 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_453
timestamp 1681620392
transform 1 0 428 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_404
timestamp 1681620392
transform 1 0 404 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_421
timestamp 1681620392
transform 1 0 388 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_294
timestamp 1681620392
transform 1 0 452 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_339
timestamp 1681620392
transform 1 0 444 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_454
timestamp 1681620392
transform 1 0 452 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_527
timestamp 1681620392
transform 1 0 444 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_552
timestamp 1681620392
transform 1 0 444 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_405
timestamp 1681620392
transform 1 0 452 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_385
timestamp 1681620392
transform 1 0 476 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_363
timestamp 1681620392
transform 1 0 476 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_455
timestamp 1681620392
transform 1 0 484 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_528
timestamp 1681620392
transform 1 0 492 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_406
timestamp 1681620392
transform 1 0 492 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_422
timestamp 1681620392
transform 1 0 492 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_295
timestamp 1681620392
transform 1 0 516 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_456
timestamp 1681620392
transform 1 0 524 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_529
timestamp 1681620392
transform 1 0 524 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_434
timestamp 1681620392
transform 1 0 508 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_296
timestamp 1681620392
transform 1 0 540 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_386
timestamp 1681620392
transform 1 0 532 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_387
timestamp 1681620392
transform 1 0 540 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_388
timestamp 1681620392
transform 1 0 556 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_340
timestamp 1681620392
transform 1 0 564 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_389
timestamp 1681620392
transform 1 0 572 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_341
timestamp 1681620392
transform 1 0 580 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_364
timestamp 1681620392
transform 1 0 556 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_384
timestamp 1681620392
transform 1 0 564 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_407
timestamp 1681620392
transform 1 0 556 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_457
timestamp 1681620392
transform 1 0 580 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_458
timestamp 1681620392
transform 1 0 588 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_530
timestamp 1681620392
transform 1 0 604 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_390
timestamp 1681620392
transform 1 0 612 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_342
timestamp 1681620392
transform 1 0 620 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_459
timestamp 1681620392
transform 1 0 612 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_460
timestamp 1681620392
transform 1 0 620 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1681620392
transform 1 0 636 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_461
timestamp 1681620392
transform 1 0 636 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_391
timestamp 1681620392
transform 1 0 660 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1681620392
transform 1 0 668 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_343
timestamp 1681620392
transform 1 0 684 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_308
timestamp 1681620392
transform 1 0 724 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_309
timestamp 1681620392
transform 1 0 740 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_310
timestamp 1681620392
transform 1 0 756 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_393
timestamp 1681620392
transform 1 0 692 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_394
timestamp 1681620392
transform 1 0 708 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_462
timestamp 1681620392
transform 1 0 684 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_531
timestamp 1681620392
transform 1 0 668 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_408
timestamp 1681620392
transform 1 0 660 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_409
timestamp 1681620392
transform 1 0 684 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_311
timestamp 1681620392
transform 1 0 812 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_395
timestamp 1681620392
transform 1 0 812 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_365
timestamp 1681620392
transform 1 0 708 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_463
timestamp 1681620392
transform 1 0 756 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_464
timestamp 1681620392
transform 1 0 788 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_366
timestamp 1681620392
transform 1 0 796 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_367
timestamp 1681620392
transform 1 0 812 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_410
timestamp 1681620392
transform 1 0 772 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_423
timestamp 1681620392
transform 1 0 724 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_424
timestamp 1681620392
transform 1 0 740 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_532
timestamp 1681620392
transform 1 0 812 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1681620392
transform 1 0 844 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_465
timestamp 1681620392
transform 1 0 844 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_368
timestamp 1681620392
transform 1 0 852 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_312
timestamp 1681620392
transform 1 0 884 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_397
timestamp 1681620392
transform 1 0 868 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_398
timestamp 1681620392
transform 1 0 884 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_344
timestamp 1681620392
transform 1 0 948 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_399
timestamp 1681620392
transform 1 0 972 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_400
timestamp 1681620392
transform 1 0 988 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_466
timestamp 1681620392
transform 1 0 860 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_467
timestamp 1681620392
transform 1 0 868 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1681620392
transform 1 0 892 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_469
timestamp 1681620392
transform 1 0 948 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_533
timestamp 1681620392
transform 1 0 852 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_411
timestamp 1681620392
transform 1 0 844 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_412
timestamp 1681620392
transform 1 0 868 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_313
timestamp 1681620392
transform 1 0 1012 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_314
timestamp 1681620392
transform 1 0 1068 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_345
timestamp 1681620392
transform 1 0 1020 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_315
timestamp 1681620392
transform 1 0 1132 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_401
timestamp 1681620392
transform 1 0 1092 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_402
timestamp 1681620392
transform 1 0 1108 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_470
timestamp 1681620392
transform 1 0 1004 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_471
timestamp 1681620392
transform 1 0 1012 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_472
timestamp 1681620392
transform 1 0 1068 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_534
timestamp 1681620392
transform 1 0 1004 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_346
timestamp 1681620392
transform 1 0 1124 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_403
timestamp 1681620392
transform 1 0 1132 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_347
timestamp 1681620392
transform 1 0 1140 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_404
timestamp 1681620392
transform 1 0 1148 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_473
timestamp 1681620392
transform 1 0 1116 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_474
timestamp 1681620392
transform 1 0 1140 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_369
timestamp 1681620392
transform 1 0 1148 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_475
timestamp 1681620392
transform 1 0 1156 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_370
timestamp 1681620392
transform 1 0 1164 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_535
timestamp 1681620392
transform 1 0 1132 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_297
timestamp 1681620392
transform 1 0 1188 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_405
timestamp 1681620392
transform 1 0 1188 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_406
timestamp 1681620392
transform 1 0 1196 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_476
timestamp 1681620392
transform 1 0 1180 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_277
timestamp 1681620392
transform 1 0 1236 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_278
timestamp 1681620392
transform 1 0 1252 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_316
timestamp 1681620392
transform 1 0 1236 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_407
timestamp 1681620392
transform 1 0 1236 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_408
timestamp 1681620392
transform 1 0 1252 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_298
timestamp 1681620392
transform 1 0 1268 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_374
timestamp 1681620392
transform 1 0 1268 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1681620392
transform 1 0 1204 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_478
timestamp 1681620392
transform 1 0 1220 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_479
timestamp 1681620392
transform 1 0 1244 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_480
timestamp 1681620392
transform 1 0 1260 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_348
timestamp 1681620392
transform 1 0 1292 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_409
timestamp 1681620392
transform 1 0 1300 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_481
timestamp 1681620392
transform 1 0 1284 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_375
timestamp 1681620392
transform 1 0 1340 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_410
timestamp 1681620392
transform 1 0 1324 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1681620392
transform 1 0 1316 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_411
timestamp 1681620392
transform 1 0 1356 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_412
timestamp 1681620392
transform 1 0 1380 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_483
timestamp 1681620392
transform 1 0 1372 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_425
timestamp 1681620392
transform 1 0 1388 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_413
timestamp 1681620392
transform 1 0 1404 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1681620392
transform 1 0 1492 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_484
timestamp 1681620392
transform 1 0 1452 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_485
timestamp 1681620392
transform 1 0 1484 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_371
timestamp 1681620392
transform 1 0 1492 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_536
timestamp 1681620392
transform 1 0 1492 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_426
timestamp 1681620392
transform 1 0 1420 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_415
timestamp 1681620392
transform 1 0 1516 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_279
timestamp 1681620392
transform 1 0 1532 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_416
timestamp 1681620392
transform 1 0 1532 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_372
timestamp 1681620392
transform 1 0 1524 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_280
timestamp 1681620392
transform 1 0 1580 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_417
timestamp 1681620392
transform 1 0 1556 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_418
timestamp 1681620392
transform 1 0 1572 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_486
timestamp 1681620392
transform 1 0 1548 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_385
timestamp 1681620392
transform 1 0 1540 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_349
timestamp 1681620392
transform 1 0 1668 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_487
timestamp 1681620392
transform 1 0 1596 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_488
timestamp 1681620392
transform 1 0 1660 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_489
timestamp 1681620392
transform 1 0 1668 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_490
timestamp 1681620392
transform 1 0 1684 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_386
timestamp 1681620392
transform 1 0 1660 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_537
timestamp 1681620392
transform 1 0 1676 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_427
timestamp 1681620392
transform 1 0 1644 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_491
timestamp 1681620392
transform 1 0 1716 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_538
timestamp 1681620392
transform 1 0 1700 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_539
timestamp 1681620392
transform 1 0 1708 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_553
timestamp 1681620392
transform 1 0 1684 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_387
timestamp 1681620392
transform 1 0 1716 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_350
timestamp 1681620392
transform 1 0 1772 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_492
timestamp 1681620392
transform 1 0 1748 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_373
timestamp 1681620392
transform 1 0 1764 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_317
timestamp 1681620392
transform 1 0 1804 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_419
timestamp 1681620392
transform 1 0 1804 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_493
timestamp 1681620392
transform 1 0 1780 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_540
timestamp 1681620392
transform 1 0 1732 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_541
timestamp 1681620392
transform 1 0 1740 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_554
timestamp 1681620392
transform 1 0 1716 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_428
timestamp 1681620392
transform 1 0 1684 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_429
timestamp 1681620392
transform 1 0 1700 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1681620392
transform 1 0 1748 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_542
timestamp 1681620392
transform 1 0 1764 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_543
timestamp 1681620392
transform 1 0 1772 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_389
timestamp 1681620392
transform 1 0 1780 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_544
timestamp 1681620392
transform 1 0 1796 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_555
timestamp 1681620392
transform 1 0 1756 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_556
timestamp 1681620392
transform 1 0 1772 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_299
timestamp 1681620392
transform 1 0 1908 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_300
timestamp 1681620392
transform 1 0 1924 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_318
timestamp 1681620392
transform 1 0 1836 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_319
timestamp 1681620392
transform 1 0 1932 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_420
timestamp 1681620392
transform 1 0 1836 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_351
timestamp 1681620392
transform 1 0 1884 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_352
timestamp 1681620392
transform 1 0 1916 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_421
timestamp 1681620392
transform 1 0 1932 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_353
timestamp 1681620392
transform 1 0 1972 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_301
timestamp 1681620392
transform 1 0 2036 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_302
timestamp 1681620392
transform 1 0 2076 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_320
timestamp 1681620392
transform 1 0 2044 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_354
timestamp 1681620392
transform 1 0 2028 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_422
timestamp 1681620392
transform 1 0 2044 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_494
timestamp 1681620392
transform 1 0 1820 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_495
timestamp 1681620392
transform 1 0 1884 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_496
timestamp 1681620392
transform 1 0 1916 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_497
timestamp 1681620392
transform 1 0 1956 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_498
timestamp 1681620392
transform 1 0 2012 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_435
timestamp 1681620392
transform 1 0 1892 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_374
timestamp 1681620392
transform 1 0 2020 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_499
timestamp 1681620392
transform 1 0 2028 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_375
timestamp 1681620392
transform 1 0 2044 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_321
timestamp 1681620392
transform 1 0 2140 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_423
timestamp 1681620392
transform 1 0 2140 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_322
timestamp 1681620392
transform 1 0 2284 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_323
timestamp 1681620392
transform 1 0 2324 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_424
timestamp 1681620392
transform 1 0 2236 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_425
timestamp 1681620392
transform 1 0 2324 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_500
timestamp 1681620392
transform 1 0 2068 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_501
timestamp 1681620392
transform 1 0 2124 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_502
timestamp 1681620392
transform 1 0 2172 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_503
timestamp 1681620392
transform 1 0 2220 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_430
timestamp 1681620392
transform 1 0 2204 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_376
timestamp 1681620392
transform 1 0 2236 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_504
timestamp 1681620392
transform 1 0 2284 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_505
timestamp 1681620392
transform 1 0 2316 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_281
timestamp 1681620392
transform 1 0 2436 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_282
timestamp 1681620392
transform 1 0 2460 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_324
timestamp 1681620392
transform 1 0 2380 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_426
timestamp 1681620392
transform 1 0 2356 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_506
timestamp 1681620392
transform 1 0 2340 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_427
timestamp 1681620392
transform 1 0 2380 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_428
timestamp 1681620392
transform 1 0 2468 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_355
timestamp 1681620392
transform 1 0 2484 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_283
timestamp 1681620392
transform 1 0 2556 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_303
timestamp 1681620392
transform 1 0 2540 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_325
timestamp 1681620392
transform 1 0 2508 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_429
timestamp 1681620392
transform 1 0 2492 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_430
timestamp 1681620392
transform 1 0 2508 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_507
timestamp 1681620392
transform 1 0 2364 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_377
timestamp 1681620392
transform 1 0 2380 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_508
timestamp 1681620392
transform 1 0 2404 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_509
timestamp 1681620392
transform 1 0 2460 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_378
timestamp 1681620392
transform 1 0 2468 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_510
timestamp 1681620392
transform 1 0 2484 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_390
timestamp 1681620392
transform 1 0 2276 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_391
timestamp 1681620392
transform 1 0 2316 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_545
timestamp 1681620392
transform 1 0 2324 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_392
timestamp 1681620392
transform 1 0 2340 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_393
timestamp 1681620392
transform 1 0 2356 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_413
timestamp 1681620392
transform 1 0 2316 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_414
timestamp 1681620392
transform 1 0 2332 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1681620392
transform 1 0 2260 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_437
timestamp 1681620392
transform 1 0 2308 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_431
timestamp 1681620392
transform 1 0 2372 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_546
timestamp 1681620392
transform 1 0 2468 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_356
timestamp 1681620392
transform 1 0 2540 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_431
timestamp 1681620392
transform 1 0 2596 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_511
timestamp 1681620392
transform 1 0 2532 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_379
timestamp 1681620392
transform 1 0 2540 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_304
timestamp 1681620392
transform 1 0 2628 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_284
timestamp 1681620392
transform 1 0 2668 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_326
timestamp 1681620392
transform 1 0 2636 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_327
timestamp 1681620392
transform 1 0 2676 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_328
timestamp 1681620392
transform 1 0 2716 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_432
timestamp 1681620392
transform 1 0 2612 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_357
timestamp 1681620392
transform 1 0 2620 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_433
timestamp 1681620392
transform 1 0 2636 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_434
timestamp 1681620392
transform 1 0 2652 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_512
timestamp 1681620392
transform 1 0 2588 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_513
timestamp 1681620392
transform 1 0 2604 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_394
timestamp 1681620392
transform 1 0 2492 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_415
timestamp 1681620392
transform 1 0 2484 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_416
timestamp 1681620392
transform 1 0 2508 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_514
timestamp 1681620392
transform 1 0 2628 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_395
timestamp 1681620392
transform 1 0 2604 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_547
timestamp 1681620392
transform 1 0 2612 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_438
timestamp 1681620392
transform 1 0 2588 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_358
timestamp 1681620392
transform 1 0 2676 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_285
timestamp 1681620392
transform 1 0 2836 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_329
timestamp 1681620392
transform 1 0 2836 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_435
timestamp 1681620392
transform 1 0 2748 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_436
timestamp 1681620392
transform 1 0 2836 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_515
timestamp 1681620392
transform 1 0 2676 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_516
timestamp 1681620392
transform 1 0 2732 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_517
timestamp 1681620392
transform 1 0 2772 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_518
timestamp 1681620392
transform 1 0 2828 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_519
timestamp 1681620392
transform 1 0 2836 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_417
timestamp 1681620392
transform 1 0 2652 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_439
timestamp 1681620392
transform 1 0 2644 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_330
timestamp 1681620392
transform 1 0 2868 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_331
timestamp 1681620392
transform 1 0 2900 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_437
timestamp 1681620392
transform 1 0 2860 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_438
timestamp 1681620392
transform 1 0 2868 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_380
timestamp 1681620392
transform 1 0 2860 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_520
timestamp 1681620392
transform 1 0 2868 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_381
timestamp 1681620392
transform 1 0 2884 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_396
timestamp 1681620392
transform 1 0 2852 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_548
timestamp 1681620392
transform 1 0 2860 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_432
timestamp 1681620392
transform 1 0 2836 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_332
timestamp 1681620392
transform 1 0 2956 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_439
timestamp 1681620392
transform 1 0 2900 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_440
timestamp 1681620392
transform 1 0 2916 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_441
timestamp 1681620392
transform 1 0 2932 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_359
timestamp 1681620392
transform 1 0 3012 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_521
timestamp 1681620392
transform 1 0 2956 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_522
timestamp 1681620392
transform 1 0 3012 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_549
timestamp 1681620392
transform 1 0 2900 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_397
timestamp 1681620392
transform 1 0 2916 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_398
timestamp 1681620392
transform 1 0 3012 0 1 2715
box -3 -3 3 3
use Project_Top_VIA0  Project_Top_VIA0_6
timestamp 1681620392
transform 1 0 24 0 1 2670
box -10 -3 10 3
use FILL  FILL_50
timestamp 1681620392
transform 1 0 72 0 -1 2770
box -8 -3 16 105
use FILL  FILL_52
timestamp 1681620392
transform 1 0 80 0 -1 2770
box -8 -3 16 105
use FILL  FILL_54
timestamp 1681620392
transform 1 0 88 0 -1 2770
box -8 -3 16 105
use FILL  FILL_56
timestamp 1681620392
transform 1 0 96 0 -1 2770
box -8 -3 16 105
use FILL  FILL_58
timestamp 1681620392
transform 1 0 104 0 -1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_9
timestamp 1681620392
transform 1 0 112 0 -1 2770
box -8 -3 40 105
use NOR2X1  NOR2X1_4
timestamp 1681620392
transform -1 0 168 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_5
timestamp 1681620392
transform -1 0 192 0 -1 2770
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_18
timestamp 1681620392
transform -1 0 288 0 -1 2770
box -8 -3 104 105
use NAND3X1  NAND3X1_10
timestamp 1681620392
transform 1 0 288 0 -1 2770
box -8 -3 40 105
use NOR2X1  NOR2X1_6
timestamp 1681620392
transform 1 0 320 0 -1 2770
box -8 -3 32 105
use INVX2  INVX2_19
timestamp 1681620392
transform 1 0 344 0 -1 2770
box -9 -3 26 105
use OAI22X1  OAI22X1_1
timestamp 1681620392
transform 1 0 360 0 -1 2770
box -8 -3 46 105
use M3_M2  M3_M2_440
timestamp 1681620392
transform 1 0 412 0 1 2675
box -3 -3 3 3
use AOI21X1  AOI21X1_1
timestamp 1681620392
transform 1 0 400 0 -1 2770
box -7 -3 39 105
use M3_M2  M3_M2_441
timestamp 1681620392
transform 1 0 444 0 1 2675
box -3 -3 3 3
use FILL  FILL_90
timestamp 1681620392
transform 1 0 432 0 -1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_11
timestamp 1681620392
transform 1 0 440 0 -1 2770
box -8 -3 40 105
use FILL  FILL_91
timestamp 1681620392
transform 1 0 472 0 -1 2770
box -8 -3 16 105
use FILL  FILL_92
timestamp 1681620392
transform 1 0 480 0 -1 2770
box -8 -3 16 105
use FILL  FILL_93
timestamp 1681620392
transform 1 0 488 0 -1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_17
timestamp 1681620392
transform 1 0 496 0 -1 2770
box -8 -3 34 105
use FILL  FILL_94
timestamp 1681620392
transform 1 0 528 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_20
timestamp 1681620392
transform 1 0 536 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_21
timestamp 1681620392
transform 1 0 552 0 -1 2770
box -9 -3 26 105
use FILL  FILL_95
timestamp 1681620392
transform 1 0 568 0 -1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_18
timestamp 1681620392
transform 1 0 576 0 -1 2770
box -8 -3 34 105
use FILL  FILL_96
timestamp 1681620392
transform 1 0 608 0 -1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_7
timestamp 1681620392
transform -1 0 640 0 -1 2770
box -8 -3 32 105
use FILL  FILL_97
timestamp 1681620392
transform 1 0 640 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_22
timestamp 1681620392
transform -1 0 664 0 -1 2770
box -9 -3 26 105
use OAI21X1  OAI21X1_19
timestamp 1681620392
transform -1 0 696 0 -1 2770
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_19
timestamp 1681620392
transform 1 0 696 0 -1 2770
box -8 -3 104 105
use NAND2X1  NAND2X1_10
timestamp 1681620392
transform 1 0 792 0 -1 2770
box -8 -3 32 105
use OAI21X1  OAI21X1_20
timestamp 1681620392
transform -1 0 848 0 -1 2770
box -8 -3 34 105
use NAND2X1  NAND2X1_11
timestamp 1681620392
transform -1 0 872 0 -1 2770
box -8 -3 32 105
use INVX2  INVX2_23
timestamp 1681620392
transform -1 0 888 0 -1 2770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_20
timestamp 1681620392
transform -1 0 984 0 -1 2770
box -8 -3 104 105
use NAND2X1  NAND2X1_12
timestamp 1681620392
transform 1 0 984 0 -1 2770
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_21
timestamp 1681620392
transform -1 0 1104 0 -1 2770
box -8 -3 104 105
use OAI21X1  OAI21X1_21
timestamp 1681620392
transform 1 0 1104 0 -1 2770
box -8 -3 34 105
use AOI22X1  AOI22X1_4
timestamp 1681620392
transform -1 0 1176 0 -1 2770
box -8 -3 46 105
use FILL  FILL_98
timestamp 1681620392
transform 1 0 1176 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_5
timestamp 1681620392
transform -1 0 1224 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_6
timestamp 1681620392
transform 1 0 1224 0 -1 2770
box -8 -3 46 105
use FILL  FILL_99
timestamp 1681620392
transform 1 0 1264 0 -1 2770
box -8 -3 16 105
use FILL  FILL_104
timestamp 1681620392
transform 1 0 1272 0 -1 2770
box -8 -3 16 105
use AOI21X1  AOI21X1_2
timestamp 1681620392
transform -1 0 1312 0 -1 2770
box -7 -3 39 105
use AOI21X1  AOI21X1_3
timestamp 1681620392
transform 1 0 1312 0 -1 2770
box -7 -3 39 105
use FILL  FILL_105
timestamp 1681620392
transform 1 0 1344 0 -1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_23
timestamp 1681620392
transform -1 0 1384 0 -1 2770
box -8 -3 34 105
use FILL  FILL_106
timestamp 1681620392
transform 1 0 1384 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_442
timestamp 1681620392
transform 1 0 1404 0 1 2675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_23
timestamp 1681620392
transform 1 0 1392 0 -1 2770
box -8 -3 104 105
use OAI21X1  OAI21X1_24
timestamp 1681620392
transform -1 0 1520 0 -1 2770
box -8 -3 34 105
use FILL  FILL_110
timestamp 1681620392
transform 1 0 1520 0 -1 2770
box -8 -3 16 105
use FILL  FILL_111
timestamp 1681620392
transform 1 0 1528 0 -1 2770
box -8 -3 16 105
use FILL  FILL_129
timestamp 1681620392
transform 1 0 1536 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_31
timestamp 1681620392
transform -1 0 1560 0 -1 2770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1681620392
transform 1 0 1560 0 -1 2770
box -8 -3 104 105
use INVX2  INVX2_32
timestamp 1681620392
transform 1 0 1656 0 -1 2770
box -9 -3 26 105
use NAND3X1  NAND3X1_12
timestamp 1681620392
transform 1 0 1672 0 -1 2770
box -8 -3 40 105
use M3_M2  M3_M2_443
timestamp 1681620392
transform 1 0 1716 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1681620392
transform 1 0 1740 0 1 2675
box -3 -3 3 3
use NAND3X1  NAND3X1_13
timestamp 1681620392
transform 1 0 1704 0 -1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_14
timestamp 1681620392
transform 1 0 1736 0 -1 2770
box -8 -3 40 105
use M3_M2  M3_M2_445
timestamp 1681620392
transform 1 0 1780 0 1 2675
box -3 -3 3 3
use NAND3X1  NAND3X1_15
timestamp 1681620392
transform 1 0 1768 0 -1 2770
box -8 -3 40 105
use BUFX2  BUFX2_0
timestamp 1681620392
transform -1 0 1824 0 -1 2770
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1681620392
transform 1 0 1824 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_31
timestamp 1681620392
transform 1 0 1920 0 -1 2770
box -8 -3 104 105
use INVX2  INVX2_33
timestamp 1681620392
transform 1 0 2016 0 -1 2770
box -9 -3 26 105
use M3_M2  M3_M2_446
timestamp 1681620392
transform 1 0 2084 0 1 2675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_32
timestamp 1681620392
transform 1 0 2032 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_33
timestamp 1681620392
transform 1 0 2128 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_34
timestamp 1681620392
transform 1 0 2224 0 -1 2770
box -8 -3 104 105
use OAI21X1  OAI21X1_39
timestamp 1681620392
transform -1 0 2352 0 -1 2770
box -8 -3 34 105
use INVX2  INVX2_34
timestamp 1681620392
transform 1 0 2352 0 -1 2770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_35
timestamp 1681620392
transform 1 0 2368 0 -1 2770
box -8 -3 104 105
use OAI21X1  OAI21X1_40
timestamp 1681620392
transform -1 0 2496 0 -1 2770
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_36
timestamp 1681620392
transform 1 0 2496 0 -1 2770
box -8 -3 104 105
use INVX2  INVX2_35
timestamp 1681620392
transform 1 0 2592 0 -1 2770
box -9 -3 26 105
use OAI21X1  OAI21X1_41
timestamp 1681620392
transform -1 0 2640 0 -1 2770
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1681620392
transform 1 0 2640 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_38
timestamp 1681620392
transform 1 0 2736 0 -1 2770
box -8 -3 104 105
use OAI21X1  OAI21X1_42
timestamp 1681620392
transform 1 0 2832 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_43
timestamp 1681620392
transform 1 0 2864 0 -1 2770
box -8 -3 34 105
use NAND2X1  NAND2X1_27
timestamp 1681620392
transform -1 0 2920 0 -1 2770
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_39
timestamp 1681620392
transform 1 0 2920 0 -1 2770
box -8 -3 104 105
use Project_Top_VIA0  Project_Top_VIA0_7
timestamp 1681620392
transform 1 0 3067 0 1 2670
box -10 -3 10 3
use M3_M2  M3_M2_501
timestamp 1681620392
transform 1 0 180 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_502
timestamp 1681620392
transform 1 0 212 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_584
timestamp 1681620392
transform 1 0 132 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_585
timestamp 1681620392
transform 1 0 172 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_586
timestamp 1681620392
transform 1 0 180 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_587
timestamp 1681620392
transform 1 0 196 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_588
timestamp 1681620392
transform 1 0 212 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_683
timestamp 1681620392
transform 1 0 84 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_562
timestamp 1681620392
transform 1 0 132 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_589
timestamp 1681620392
transform 1 0 236 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1681620392
transform 1 0 252 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_447
timestamp 1681620392
transform 1 0 276 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_503
timestamp 1681620392
transform 1 0 276 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_504
timestamp 1681620392
transform 1 0 300 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_591
timestamp 1681620392
transform 1 0 276 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1681620392
transform 1 0 308 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_684
timestamp 1681620392
transform 1 0 188 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_685
timestamp 1681620392
transform 1 0 204 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_686
timestamp 1681620392
transform 1 0 220 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_687
timestamp 1681620392
transform 1 0 228 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_688
timestamp 1681620392
transform 1 0 244 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1681620392
transform 1 0 268 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1681620392
transform 1 0 284 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_691
timestamp 1681620392
transform 1 0 300 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_563
timestamp 1681620392
transform 1 0 204 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_564
timestamp 1681620392
transform 1 0 220 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_598
timestamp 1681620392
transform 1 0 188 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_565
timestamp 1681620392
transform 1 0 268 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_599
timestamp 1681620392
transform 1 0 228 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_600
timestamp 1681620392
transform 1 0 300 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_525
timestamp 1681620392
transform 1 0 316 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_464
timestamp 1681620392
transform 1 0 356 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_593
timestamp 1681620392
transform 1 0 324 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1681620392
transform 1 0 340 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1681620392
transform 1 0 348 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_692
timestamp 1681620392
transform 1 0 316 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_693
timestamp 1681620392
transform 1 0 332 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_545
timestamp 1681620392
transform 1 0 340 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_694
timestamp 1681620392
transform 1 0 348 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_546
timestamp 1681620392
transform 1 0 356 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_566
timestamp 1681620392
transform 1 0 348 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_596
timestamp 1681620392
transform 1 0 372 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_778
timestamp 1681620392
transform 1 0 380 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_505
timestamp 1681620392
transform 1 0 404 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_695
timestamp 1681620392
transform 1 0 404 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_506
timestamp 1681620392
transform 1 0 444 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_597
timestamp 1681620392
transform 1 0 436 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_598
timestamp 1681620392
transform 1 0 444 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_696
timestamp 1681620392
transform 1 0 428 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_779
timestamp 1681620392
transform 1 0 412 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_567
timestamp 1681620392
transform 1 0 420 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_601
timestamp 1681620392
transform 1 0 412 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_697
timestamp 1681620392
transform 1 0 452 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_599
timestamp 1681620392
transform 1 0 476 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_780
timestamp 1681620392
transform 1 0 468 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_602
timestamp 1681620392
transform 1 0 468 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_698
timestamp 1681620392
transform 1 0 492 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_557
timestamp 1681620392
transform 1 0 532 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_558
timestamp 1681620392
transform 1 0 548 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_559
timestamp 1681620392
transform 1 0 516 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_560
timestamp 1681620392
transform 1 0 540 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_561
timestamp 1681620392
transform 1 0 556 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_600
timestamp 1681620392
transform 1 0 508 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1681620392
transform 1 0 524 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_526
timestamp 1681620392
transform 1 0 532 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_602
timestamp 1681620392
transform 1 0 556 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_562
timestamp 1681620392
transform 1 0 580 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_568
timestamp 1681620392
transform 1 0 580 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_603
timestamp 1681620392
transform 1 0 588 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_478
timestamp 1681620392
transform 1 0 620 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_479
timestamp 1681620392
transform 1 0 636 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_563
timestamp 1681620392
transform 1 0 652 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_604
timestamp 1681620392
transform 1 0 620 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_605
timestamp 1681620392
transform 1 0 636 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_699
timestamp 1681620392
transform 1 0 612 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_700
timestamp 1681620392
transform 1 0 628 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_781
timestamp 1681620392
transform 1 0 596 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_603
timestamp 1681620392
transform 1 0 596 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_569
timestamp 1681620392
transform 1 0 628 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_701
timestamp 1681620392
transform 1 0 652 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_604
timestamp 1681620392
transform 1 0 644 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_480
timestamp 1681620392
transform 1 0 668 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_782
timestamp 1681620392
transform 1 0 668 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_606
timestamp 1681620392
transform 1 0 692 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_702
timestamp 1681620392
transform 1 0 700 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_465
timestamp 1681620392
transform 1 0 756 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_607
timestamp 1681620392
transform 1 0 716 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_527
timestamp 1681620392
transform 1 0 724 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_608
timestamp 1681620392
transform 1 0 772 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_703
timestamp 1681620392
transform 1 0 796 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_570
timestamp 1681620392
transform 1 0 772 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_564
timestamp 1681620392
transform 1 0 836 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_528
timestamp 1681620392
transform 1 0 820 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_704
timestamp 1681620392
transform 1 0 820 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_705
timestamp 1681620392
transform 1 0 836 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_448
timestamp 1681620392
transform 1 0 860 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_449
timestamp 1681620392
transform 1 0 972 0 1 2665
box -3 -3 3 3
use M2_M1  M2_M1_565
timestamp 1681620392
transform 1 0 972 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_609
timestamp 1681620392
transform 1 0 860 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1681620392
transform 1 0 876 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1681620392
transform 1 0 932 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_571
timestamp 1681620392
transform 1 0 836 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_706
timestamp 1681620392
transform 1 0 868 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_707
timestamp 1681620392
transform 1 0 956 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_708
timestamp 1681620392
transform 1 0 972 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_605
timestamp 1681620392
transform 1 0 860 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_572
timestamp 1681620392
transform 1 0 932 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_573
timestamp 1681620392
transform 1 0 972 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_612
timestamp 1681620392
transform 1 0 1004 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_709
timestamp 1681620392
transform 1 0 996 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_547
timestamp 1681620392
transform 1 0 1004 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_529
timestamp 1681620392
transform 1 0 1020 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_613
timestamp 1681620392
transform 1 0 1068 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_530
timestamp 1681620392
transform 1 0 1092 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_614
timestamp 1681620392
transform 1 0 1108 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_615
timestamp 1681620392
transform 1 0 1116 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_616
timestamp 1681620392
transform 1 0 1124 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_710
timestamp 1681620392
transform 1 0 1020 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_574
timestamp 1681620392
transform 1 0 1068 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_548
timestamp 1681620392
transform 1 0 1116 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_481
timestamp 1681620392
transform 1 0 1156 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_507
timestamp 1681620392
transform 1 0 1148 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_531
timestamp 1681620392
transform 1 0 1140 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_508
timestamp 1681620392
transform 1 0 1188 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_566
timestamp 1681620392
transform 1 0 1204 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_617
timestamp 1681620392
transform 1 0 1156 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_532
timestamp 1681620392
transform 1 0 1180 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_618
timestamp 1681620392
transform 1 0 1188 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_619
timestamp 1681620392
transform 1 0 1204 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_711
timestamp 1681620392
transform 1 0 1140 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_712
timestamp 1681620392
transform 1 0 1148 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_549
timestamp 1681620392
transform 1 0 1156 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_713
timestamp 1681620392
transform 1 0 1172 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_714
timestamp 1681620392
transform 1 0 1180 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_715
timestamp 1681620392
transform 1 0 1204 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_783
timestamp 1681620392
transform 1 0 1140 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_575
timestamp 1681620392
transform 1 0 1204 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_482
timestamp 1681620392
transform 1 0 1220 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_620
timestamp 1681620392
transform 1 0 1220 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_621
timestamp 1681620392
transform 1 0 1244 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_716
timestamp 1681620392
transform 1 0 1228 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_717
timestamp 1681620392
transform 1 0 1236 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_576
timestamp 1681620392
transform 1 0 1228 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_550
timestamp 1681620392
transform 1 0 1244 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_450
timestamp 1681620392
transform 1 0 1284 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_454
timestamp 1681620392
transform 1 0 1276 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_466
timestamp 1681620392
transform 1 0 1268 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_467
timestamp 1681620392
transform 1 0 1300 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_483
timestamp 1681620392
transform 1 0 1268 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_718
timestamp 1681620392
transform 1 0 1260 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_606
timestamp 1681620392
transform 1 0 1236 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_577
timestamp 1681620392
transform 1 0 1260 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_567
timestamp 1681620392
transform 1 0 1268 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_622
timestamp 1681620392
transform 1 0 1268 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_623
timestamp 1681620392
transform 1 0 1292 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_719
timestamp 1681620392
transform 1 0 1276 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_607
timestamp 1681620392
transform 1 0 1268 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_484
timestamp 1681620392
transform 1 0 1308 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_624
timestamp 1681620392
transform 1 0 1308 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_720
timestamp 1681620392
transform 1 0 1300 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_551
timestamp 1681620392
transform 1 0 1308 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_721
timestamp 1681620392
transform 1 0 1316 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_784
timestamp 1681620392
transform 1 0 1308 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_608
timestamp 1681620392
transform 1 0 1316 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_451
timestamp 1681620392
transform 1 0 1340 0 1 2665
box -3 -3 3 3
use M2_M1  M2_M1_568
timestamp 1681620392
transform 1 0 1340 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_485
timestamp 1681620392
transform 1 0 1356 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_569
timestamp 1681620392
transform 1 0 1348 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_625
timestamp 1681620392
transform 1 0 1356 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_722
timestamp 1681620392
transform 1 0 1340 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_552
timestamp 1681620392
transform 1 0 1348 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_455
timestamp 1681620392
transform 1 0 1388 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_570
timestamp 1681620392
transform 1 0 1388 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_626
timestamp 1681620392
transform 1 0 1380 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_723
timestamp 1681620392
transform 1 0 1380 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_578
timestamp 1681620392
transform 1 0 1380 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_627
timestamp 1681620392
transform 1 0 1412 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_724
timestamp 1681620392
transform 1 0 1404 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_579
timestamp 1681620392
transform 1 0 1404 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_725
timestamp 1681620392
transform 1 0 1420 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_571
timestamp 1681620392
transform 1 0 1436 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_509
timestamp 1681620392
transform 1 0 1444 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1681620392
transform 1 0 1436 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_533
timestamp 1681620392
transform 1 0 1452 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_510
timestamp 1681620392
transform 1 0 1484 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_572
timestamp 1681620392
transform 1 0 1492 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_534
timestamp 1681620392
transform 1 0 1492 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_726
timestamp 1681620392
transform 1 0 1476 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_727
timestamp 1681620392
transform 1 0 1492 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_728
timestamp 1681620392
transform 1 0 1524 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_628
timestamp 1681620392
transform 1 0 1540 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_468
timestamp 1681620392
transform 1 0 1556 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_573
timestamp 1681620392
transform 1 0 1572 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_629
timestamp 1681620392
transform 1 0 1556 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_729
timestamp 1681620392
transform 1 0 1548 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_610
timestamp 1681620392
transform 1 0 1540 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_469
timestamp 1681620392
transform 1 0 1668 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_535
timestamp 1681620392
transform 1 0 1588 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_630
timestamp 1681620392
transform 1 0 1612 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_631
timestamp 1681620392
transform 1 0 1668 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_632
timestamp 1681620392
transform 1 0 1676 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_730
timestamp 1681620392
transform 1 0 1572 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_731
timestamp 1681620392
transform 1 0 1588 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_580
timestamp 1681620392
transform 1 0 1572 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_581
timestamp 1681620392
transform 1 0 1612 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_470
timestamp 1681620392
transform 1 0 1772 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_471
timestamp 1681620392
transform 1 0 1820 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_472
timestamp 1681620392
transform 1 0 1844 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_486
timestamp 1681620392
transform 1 0 1804 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_511
timestamp 1681620392
transform 1 0 1732 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_512
timestamp 1681620392
transform 1 0 1788 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_536
timestamp 1681620392
transform 1 0 1700 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_633
timestamp 1681620392
transform 1 0 1724 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_634
timestamp 1681620392
transform 1 0 1780 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1681620392
transform 1 0 1788 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_732
timestamp 1681620392
transform 1 0 1684 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_733
timestamp 1681620392
transform 1 0 1700 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_582
timestamp 1681620392
transform 1 0 1684 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_553
timestamp 1681620392
transform 1 0 1780 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_734
timestamp 1681620392
transform 1 0 1788 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_611
timestamp 1681620392
transform 1 0 1724 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_612
timestamp 1681620392
transform 1 0 1772 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_574
timestamp 1681620392
transform 1 0 1812 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_513
timestamp 1681620392
transform 1 0 1820 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_537
timestamp 1681620392
transform 1 0 1812 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_636
timestamp 1681620392
transform 1 0 1828 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_637
timestamp 1681620392
transform 1 0 1876 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_538
timestamp 1681620392
transform 1 0 1892 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_638
timestamp 1681620392
transform 1 0 1924 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_639
timestamp 1681620392
transform 1 0 1932 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_735
timestamp 1681620392
transform 1 0 1812 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_736
timestamp 1681620392
transform 1 0 1820 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_583
timestamp 1681620392
transform 1 0 1796 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_554
timestamp 1681620392
transform 1 0 1828 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_737
timestamp 1681620392
transform 1 0 1844 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_487
timestamp 1681620392
transform 1 0 1948 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_488
timestamp 1681620392
transform 1 0 1964 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_575
timestamp 1681620392
transform 1 0 1948 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_456
timestamp 1681620392
transform 1 0 1988 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_457
timestamp 1681620392
transform 1 0 2012 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_514
timestamp 1681620392
transform 1 0 1980 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_489
timestamp 1681620392
transform 1 0 2036 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_576
timestamp 1681620392
transform 1 0 2020 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_640
timestamp 1681620392
transform 1 0 1964 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1681620392
transform 1 0 1980 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1681620392
transform 1 0 1996 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_643
timestamp 1681620392
transform 1 0 2012 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_738
timestamp 1681620392
transform 1 0 1940 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_739
timestamp 1681620392
transform 1 0 1948 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_584
timestamp 1681620392
transform 1 0 1908 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_585
timestamp 1681620392
transform 1 0 1924 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_586
timestamp 1681620392
transform 1 0 1940 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_613
timestamp 1681620392
transform 1 0 1828 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_539
timestamp 1681620392
transform 1 0 2020 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_644
timestamp 1681620392
transform 1 0 2036 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1681620392
transform 1 0 2044 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_740
timestamp 1681620392
transform 1 0 1972 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_555
timestamp 1681620392
transform 1 0 1980 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_741
timestamp 1681620392
transform 1 0 1988 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_556
timestamp 1681620392
transform 1 0 1996 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_742
timestamp 1681620392
transform 1 0 2004 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_743
timestamp 1681620392
transform 1 0 2020 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_614
timestamp 1681620392
transform 1 0 2036 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_452
timestamp 1681620392
transform 1 0 2092 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_490
timestamp 1681620392
transform 1 0 2060 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_491
timestamp 1681620392
transform 1 0 2076 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_458
timestamp 1681620392
transform 1 0 2108 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_515
timestamp 1681620392
transform 1 0 2076 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_516
timestamp 1681620392
transform 1 0 2100 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_540
timestamp 1681620392
transform 1 0 2068 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_459
timestamp 1681620392
transform 1 0 2156 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_492
timestamp 1681620392
transform 1 0 2116 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_646
timestamp 1681620392
transform 1 0 2076 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_647
timestamp 1681620392
transform 1 0 2092 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_648
timestamp 1681620392
transform 1 0 2108 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_744
timestamp 1681620392
transform 1 0 2076 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_745
timestamp 1681620392
transform 1 0 2084 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_746
timestamp 1681620392
transform 1 0 2100 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_517
timestamp 1681620392
transform 1 0 2124 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_493
timestamp 1681620392
transform 1 0 2164 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_577
timestamp 1681620392
transform 1 0 2164 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_649
timestamp 1681620392
transform 1 0 2140 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_650
timestamp 1681620392
transform 1 0 2156 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_651
timestamp 1681620392
transform 1 0 2180 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_652
timestamp 1681620392
transform 1 0 2188 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_653
timestamp 1681620392
transform 1 0 2204 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_747
timestamp 1681620392
transform 1 0 2124 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_748
timestamp 1681620392
transform 1 0 2156 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_749
timestamp 1681620392
transform 1 0 2164 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_785
timestamp 1681620392
transform 1 0 2116 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_587
timestamp 1681620392
transform 1 0 2124 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_588
timestamp 1681620392
transform 1 0 2156 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_750
timestamp 1681620392
transform 1 0 2204 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_589
timestamp 1681620392
transform 1 0 2204 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_615
timestamp 1681620392
transform 1 0 2180 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_473
timestamp 1681620392
transform 1 0 2236 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_751
timestamp 1681620392
transform 1 0 2220 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_752
timestamp 1681620392
transform 1 0 2228 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_578
timestamp 1681620392
transform 1 0 2260 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_654
timestamp 1681620392
transform 1 0 2244 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_655
timestamp 1681620392
transform 1 0 2260 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_753
timestamp 1681620392
transform 1 0 2260 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_460
timestamp 1681620392
transform 1 0 2300 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_494
timestamp 1681620392
transform 1 0 2284 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_579
timestamp 1681620392
transform 1 0 2308 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_656
timestamp 1681620392
transform 1 0 2284 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_657
timestamp 1681620392
transform 1 0 2292 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_557
timestamp 1681620392
transform 1 0 2276 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_754
timestamp 1681620392
transform 1 0 2284 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_616
timestamp 1681620392
transform 1 0 2284 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_474
timestamp 1681620392
transform 1 0 2332 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_461
timestamp 1681620392
transform 1 0 2372 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_495
timestamp 1681620392
transform 1 0 2356 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_518
timestamp 1681620392
transform 1 0 2324 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_519
timestamp 1681620392
transform 1 0 2364 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_658
timestamp 1681620392
transform 1 0 2332 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_659
timestamp 1681620392
transform 1 0 2348 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_660
timestamp 1681620392
transform 1 0 2364 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_661
timestamp 1681620392
transform 1 0 2372 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_755
timestamp 1681620392
transform 1 0 2308 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_756
timestamp 1681620392
transform 1 0 2316 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_617
timestamp 1681620392
transform 1 0 2308 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_757
timestamp 1681620392
transform 1 0 2340 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_558
timestamp 1681620392
transform 1 0 2348 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_496
timestamp 1681620392
transform 1 0 2388 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_580
timestamp 1681620392
transform 1 0 2388 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_581
timestamp 1681620392
transform 1 0 2420 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_662
timestamp 1681620392
transform 1 0 2404 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_758
timestamp 1681620392
transform 1 0 2372 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_559
timestamp 1681620392
transform 1 0 2380 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_759
timestamp 1681620392
transform 1 0 2388 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_475
timestamp 1681620392
transform 1 0 2436 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_520
timestamp 1681620392
transform 1 0 2436 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_497
timestamp 1681620392
transform 1 0 2476 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_663
timestamp 1681620392
transform 1 0 2428 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_664
timestamp 1681620392
transform 1 0 2436 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1681620392
transform 1 0 2460 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_666
timestamp 1681620392
transform 1 0 2476 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_760
timestamp 1681620392
transform 1 0 2412 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_590
timestamp 1681620392
transform 1 0 2420 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_618
timestamp 1681620392
transform 1 0 2404 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_761
timestamp 1681620392
transform 1 0 2444 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_762
timestamp 1681620392
transform 1 0 2452 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_763
timestamp 1681620392
transform 1 0 2484 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_462
timestamp 1681620392
transform 1 0 2492 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_476
timestamp 1681620392
transform 1 0 2556 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_453
timestamp 1681620392
transform 1 0 2604 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_477
timestamp 1681620392
transform 1 0 2612 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_521
timestamp 1681620392
transform 1 0 2596 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_498
timestamp 1681620392
transform 1 0 2628 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_499
timestamp 1681620392
transform 1 0 2668 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_500
timestamp 1681620392
transform 1 0 2708 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_522
timestamp 1681620392
transform 1 0 2636 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_523
timestamp 1681620392
transform 1 0 2660 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_524
timestamp 1681620392
transform 1 0 2676 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_667
timestamp 1681620392
transform 1 0 2492 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1681620392
transform 1 0 2540 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_669
timestamp 1681620392
transform 1 0 2588 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_670
timestamp 1681620392
transform 1 0 2596 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_671
timestamp 1681620392
transform 1 0 2612 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_672
timestamp 1681620392
transform 1 0 2628 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_673
timestamp 1681620392
transform 1 0 2636 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_674
timestamp 1681620392
transform 1 0 2652 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_675
timestamp 1681620392
transform 1 0 2668 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_676
timestamp 1681620392
transform 1 0 2676 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_764
timestamp 1681620392
transform 1 0 2508 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_765
timestamp 1681620392
transform 1 0 2596 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_766
timestamp 1681620392
transform 1 0 2620 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_591
timestamp 1681620392
transform 1 0 2596 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_592
timestamp 1681620392
transform 1 0 2620 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_541
timestamp 1681620392
transform 1 0 2684 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_677
timestamp 1681620392
transform 1 0 2692 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_678
timestamp 1681620392
transform 1 0 2708 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_679
timestamp 1681620392
transform 1 0 2716 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_767
timestamp 1681620392
transform 1 0 2644 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_768
timestamp 1681620392
transform 1 0 2676 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_769
timestamp 1681620392
transform 1 0 2684 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_770
timestamp 1681620392
transform 1 0 2700 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_593
timestamp 1681620392
transform 1 0 2676 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_582
timestamp 1681620392
transform 1 0 2732 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_771
timestamp 1681620392
transform 1 0 2724 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_560
timestamp 1681620392
transform 1 0 2740 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_680
timestamp 1681620392
transform 1 0 2780 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_542
timestamp 1681620392
transform 1 0 2796 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_772
timestamp 1681620392
transform 1 0 2764 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_561
timestamp 1681620392
transform 1 0 2780 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_773
timestamp 1681620392
transform 1 0 2796 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_594
timestamp 1681620392
transform 1 0 2796 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_595
timestamp 1681620392
transform 1 0 2828 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_774
timestamp 1681620392
transform 1 0 2844 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_463
timestamp 1681620392
transform 1 0 2868 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_583
timestamp 1681620392
transform 1 0 2876 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_775
timestamp 1681620392
transform 1 0 2876 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_596
timestamp 1681620392
transform 1 0 2876 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_543
timestamp 1681620392
transform 1 0 2916 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_776
timestamp 1681620392
transform 1 0 2916 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_681
timestamp 1681620392
transform 1 0 2956 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_544
timestamp 1681620392
transform 1 0 3004 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_682
timestamp 1681620392
transform 1 0 3012 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_777
timestamp 1681620392
transform 1 0 2932 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_597
timestamp 1681620392
transform 1 0 2956 0 1 2595
box -3 -3 3 3
use Project_Top_VIA0  Project_Top_VIA0_8
timestamp 1681620392
transform 1 0 48 0 1 2570
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_40
timestamp 1681620392
transform 1 0 72 0 1 2570
box -8 -3 104 105
use INVX2  INVX2_36
timestamp 1681620392
transform 1 0 168 0 1 2570
box -9 -3 26 105
use OAI22X1  OAI22X1_2
timestamp 1681620392
transform 1 0 184 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_3
timestamp 1681620392
transform 1 0 224 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_4
timestamp 1681620392
transform -1 0 304 0 1 2570
box -8 -3 46 105
use FILL  FILL_130
timestamp 1681620392
transform 1 0 304 0 1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_5
timestamp 1681620392
transform -1 0 352 0 1 2570
box -8 -3 46 105
use NOR2X1  NOR2X1_10
timestamp 1681620392
transform -1 0 376 0 1 2570
box -8 -3 32 105
use FILL  FILL_131
timestamp 1681620392
transform 1 0 376 0 1 2570
box -8 -3 16 105
use FILL  FILL_132
timestamp 1681620392
transform 1 0 384 0 1 2570
box -8 -3 16 105
use FILL  FILL_133
timestamp 1681620392
transform 1 0 392 0 1 2570
box -8 -3 16 105
use FILL  FILL_134
timestamp 1681620392
transform 1 0 400 0 1 2570
box -8 -3 16 105
use AOI21X1  AOI21X1_4
timestamp 1681620392
transform -1 0 440 0 1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_5
timestamp 1681620392
transform 1 0 440 0 1 2570
box -7 -3 39 105
use FILL  FILL_135
timestamp 1681620392
transform 1 0 472 0 1 2570
box -8 -3 16 105
use FILL  FILL_136
timestamp 1681620392
transform 1 0 480 0 1 2570
box -8 -3 16 105
use FILL  FILL_137
timestamp 1681620392
transform 1 0 488 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_38
timestamp 1681620392
transform 1 0 496 0 1 2570
box -9 -3 26 105
use NAND3X1  NAND3X1_16
timestamp 1681620392
transform 1 0 512 0 1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_17
timestamp 1681620392
transform 1 0 544 0 1 2570
box -8 -3 40 105
use FILL  FILL_138
timestamp 1681620392
transform 1 0 576 0 1 2570
box -8 -3 16 105
use FILL  FILL_139
timestamp 1681620392
transform 1 0 584 0 1 2570
box -8 -3 16 105
use AOI21X1  AOI21X1_6
timestamp 1681620392
transform -1 0 624 0 1 2570
box -7 -3 39 105
use OAI21X1  OAI21X1_44
timestamp 1681620392
transform 1 0 624 0 1 2570
box -8 -3 34 105
use FILL  FILL_146
timestamp 1681620392
transform 1 0 656 0 1 2570
box -8 -3 16 105
use FILL  FILL_148
timestamp 1681620392
transform 1 0 664 0 1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_11
timestamp 1681620392
transform 1 0 672 0 1 2570
box -8 -3 32 105
use FILL  FILL_149
timestamp 1681620392
transform 1 0 696 0 1 2570
box -8 -3 16 105
use FILL  FILL_150
timestamp 1681620392
transform 1 0 704 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_619
timestamp 1681620392
transform 1 0 796 0 1 2575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_45
timestamp 1681620392
transform -1 0 808 0 1 2570
box -8 -3 104 105
use FILL  FILL_153
timestamp 1681620392
transform 1 0 808 0 1 2570
box -8 -3 16 105
use NAND2X1  NAND2X1_28
timestamp 1681620392
transform 1 0 816 0 1 2570
box -8 -3 32 105
use OAI21X1  OAI21X1_47
timestamp 1681620392
transform -1 0 872 0 1 2570
box -8 -3 34 105
use M3_M2  M3_M2_620
timestamp 1681620392
transform 1 0 956 0 1 2575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_46
timestamp 1681620392
transform -1 0 968 0 1 2570
box -8 -3 104 105
use OAI21X1  OAI21X1_48
timestamp 1681620392
transform -1 0 1000 0 1 2570
box -8 -3 34 105
use FILL  FILL_154
timestamp 1681620392
transform 1 0 1000 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_621
timestamp 1681620392
transform 1 0 1044 0 1 2575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_47
timestamp 1681620392
transform 1 0 1008 0 1 2570
box -8 -3 104 105
use INVX2  INVX2_43
timestamp 1681620392
transform 1 0 1104 0 1 2570
box -9 -3 26 105
use NOR2X1  NOR2X1_13
timestamp 1681620392
transform -1 0 1144 0 1 2570
box -8 -3 32 105
use OAI21X1  OAI21X1_49
timestamp 1681620392
transform 1 0 1144 0 1 2570
box -8 -3 34 105
use M3_M2  M3_M2_622
timestamp 1681620392
transform 1 0 1196 0 1 2575
box -3 -3 3 3
use OAI21X1  OAI21X1_50
timestamp 1681620392
transform 1 0 1176 0 1 2570
box -8 -3 34 105
use INVX2  INVX2_45
timestamp 1681620392
transform -1 0 1224 0 1 2570
box -9 -3 26 105
use FILL  FILL_164
timestamp 1681620392
transform 1 0 1224 0 1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_51
timestamp 1681620392
transform 1 0 1232 0 1 2570
box -8 -3 34 105
use FILL  FILL_169
timestamp 1681620392
transform 1 0 1264 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_46
timestamp 1681620392
transform 1 0 1272 0 1 2570
box -9 -3 26 105
use NOR2X1  NOR2X1_14
timestamp 1681620392
transform -1 0 1312 0 1 2570
box -8 -3 32 105
use OAI21X1  OAI21X1_52
timestamp 1681620392
transform 1 0 1312 0 1 2570
box -8 -3 34 105
use FILL  FILL_170
timestamp 1681620392
transform 1 0 1344 0 1 2570
box -8 -3 16 105
use FILL  FILL_171
timestamp 1681620392
transform 1 0 1352 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_623
timestamp 1681620392
transform 1 0 1388 0 1 2575
box -3 -3 3 3
use NAND2X1  NAND2X1_30
timestamp 1681620392
transform -1 0 1384 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_31
timestamp 1681620392
transform -1 0 1408 0 1 2570
box -8 -3 32 105
use FILL  FILL_172
timestamp 1681620392
transform 1 0 1408 0 1 2570
box -8 -3 16 105
use NAND2X1  NAND2X1_32
timestamp 1681620392
transform 1 0 1416 0 1 2570
box -8 -3 32 105
use FILL  FILL_173
timestamp 1681620392
transform 1 0 1440 0 1 2570
box -8 -3 16 105
use FILL  FILL_181
timestamp 1681620392
transform 1 0 1448 0 1 2570
box -8 -3 16 105
use FILL  FILL_183
timestamp 1681620392
transform 1 0 1456 0 1 2570
box -8 -3 16 105
use FILL  FILL_184
timestamp 1681620392
transform 1 0 1464 0 1 2570
box -8 -3 16 105
use NAND2X1  NAND2X1_33
timestamp 1681620392
transform 1 0 1472 0 1 2570
box -8 -3 32 105
use OAI21X1  OAI21X1_54
timestamp 1681620392
transform -1 0 1528 0 1 2570
box -8 -3 34 105
use FILL  FILL_185
timestamp 1681620392
transform 1 0 1528 0 1 2570
box -8 -3 16 105
use FILL  FILL_186
timestamp 1681620392
transform 1 0 1536 0 1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_55
timestamp 1681620392
transform 1 0 1544 0 1 2570
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_51
timestamp 1681620392
transform 1 0 1576 0 1 2570
box -8 -3 104 105
use INVX2  INVX2_48
timestamp 1681620392
transform -1 0 1688 0 1 2570
box -9 -3 26 105
use M3_M2  M3_M2_624
timestamp 1681620392
transform 1 0 1788 0 1 2575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_53
timestamp 1681620392
transform 1 0 1688 0 1 2570
box -8 -3 104 105
use OAI21X1  OAI21X1_58
timestamp 1681620392
transform 1 0 1784 0 1 2570
box -8 -3 34 105
use INVX2  INVX2_49
timestamp 1681620392
transform 1 0 1816 0 1 2570
box -9 -3 26 105
use M3_M2  M3_M2_625
timestamp 1681620392
transform 1 0 1900 0 1 2575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_54
timestamp 1681620392
transform 1 0 1832 0 1 2570
box -8 -3 104 105
use INVX2  INVX2_50
timestamp 1681620392
transform -1 0 1944 0 1 2570
box -9 -3 26 105
use OAI21X1  OAI21X1_59
timestamp 1681620392
transform -1 0 1976 0 1 2570
box -8 -3 34 105
use AOI22X1  AOI22X1_7
timestamp 1681620392
transform 1 0 1976 0 1 2570
box -8 -3 46 105
use OAI21X1  OAI21X1_60
timestamp 1681620392
transform -1 0 2048 0 1 2570
box -8 -3 34 105
use FILL  FILL_189
timestamp 1681620392
transform 1 0 2048 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_51
timestamp 1681620392
transform -1 0 2072 0 1 2570
box -9 -3 26 105
use AOI22X1  AOI22X1_8
timestamp 1681620392
transform 1 0 2072 0 1 2570
box -8 -3 46 105
use FILL  FILL_190
timestamp 1681620392
transform 1 0 2112 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_9
timestamp 1681620392
transform 1 0 2120 0 1 2570
box -8 -3 46 105
use OAI21X1  OAI21X1_61
timestamp 1681620392
transform -1 0 2192 0 1 2570
box -8 -3 34 105
use INVX2  INVX2_52
timestamp 1681620392
transform -1 0 2208 0 1 2570
box -9 -3 26 105
use FILL  FILL_191
timestamp 1681620392
transform 1 0 2208 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_626
timestamp 1681620392
transform 1 0 2228 0 1 2575
box -3 -3 3 3
use FILL  FILL_192
timestamp 1681620392
transform 1 0 2216 0 1 2570
box -8 -3 16 105
use FILL  FILL_193
timestamp 1681620392
transform 1 0 2224 0 1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_62
timestamp 1681620392
transform 1 0 2232 0 1 2570
box -8 -3 34 105
use M3_M2  M3_M2_627
timestamp 1681620392
transform 1 0 2292 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_628
timestamp 1681620392
transform 1 0 2316 0 1 2575
box -3 -3 3 3
use INVX2  INVX2_53
timestamp 1681620392
transform 1 0 2264 0 1 2570
box -9 -3 26 105
use OAI21X1  OAI21X1_63
timestamp 1681620392
transform 1 0 2280 0 1 2570
box -8 -3 34 105
use INVX2  INVX2_54
timestamp 1681620392
transform 1 0 2312 0 1 2570
box -9 -3 26 105
use AOI22X1  AOI22X1_10
timestamp 1681620392
transform 1 0 2328 0 1 2570
box -8 -3 46 105
use INVX2  INVX2_55
timestamp 1681620392
transform 1 0 2368 0 1 2570
box -9 -3 26 105
use OAI21X1  OAI21X1_64
timestamp 1681620392
transform -1 0 2416 0 1 2570
box -8 -3 34 105
use NAND2X1  NAND2X1_35
timestamp 1681620392
transform -1 0 2440 0 1 2570
box -8 -3 32 105
use AOI22X1  AOI22X1_11
timestamp 1681620392
transform 1 0 2440 0 1 2570
box -8 -3 46 105
use INVX2  INVX2_56
timestamp 1681620392
transform 1 0 2480 0 1 2570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_55
timestamp 1681620392
transform 1 0 2496 0 1 2570
box -8 -3 104 105
use AOI22X1  AOI22X1_12
timestamp 1681620392
transform 1 0 2592 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_13
timestamp 1681620392
transform 1 0 2632 0 1 2570
box -8 -3 46 105
use M3_M2  M3_M2_629
timestamp 1681620392
transform 1 0 2684 0 1 2575
box -3 -3 3 3
use AOI22X1  AOI22X1_14
timestamp 1681620392
transform 1 0 2672 0 1 2570
box -8 -3 46 105
use M3_M2  M3_M2_630
timestamp 1681620392
transform 1 0 2724 0 1 2575
box -3 -3 3 3
use INVX2  INVX2_57
timestamp 1681620392
transform -1 0 2728 0 1 2570
box -9 -3 26 105
use FILL  FILL_194
timestamp 1681620392
transform 1 0 2728 0 1 2570
box -8 -3 16 105
use FILL  FILL_195
timestamp 1681620392
transform 1 0 2736 0 1 2570
box -8 -3 16 105
use FILL  FILL_196
timestamp 1681620392
transform 1 0 2744 0 1 2570
box -8 -3 16 105
use FILL  FILL_197
timestamp 1681620392
transform 1 0 2752 0 1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_65
timestamp 1681620392
transform -1 0 2792 0 1 2570
box -8 -3 34 105
use INVX2  INVX2_58
timestamp 1681620392
transform 1 0 2792 0 1 2570
box -9 -3 26 105
use FILL  FILL_198
timestamp 1681620392
transform 1 0 2808 0 1 2570
box -8 -3 16 105
use FILL  FILL_199
timestamp 1681620392
transform 1 0 2816 0 1 2570
box -8 -3 16 105
use FILL  FILL_200
timestamp 1681620392
transform 1 0 2824 0 1 2570
box -8 -3 16 105
use FILL  FILL_201
timestamp 1681620392
transform 1 0 2832 0 1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_66
timestamp 1681620392
transform 1 0 2840 0 1 2570
box -8 -3 34 105
use NAND2X1  NAND2X1_36
timestamp 1681620392
transform -1 0 2896 0 1 2570
box -8 -3 32 105
use FILL  FILL_202
timestamp 1681620392
transform 1 0 2896 0 1 2570
box -8 -3 16 105
use FILL  FILL_203
timestamp 1681620392
transform 1 0 2904 0 1 2570
box -8 -3 16 105
use FILL  FILL_204
timestamp 1681620392
transform 1 0 2912 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_56
timestamp 1681620392
transform 1 0 2920 0 1 2570
box -8 -3 104 105
use Project_Top_VIA0  Project_Top_VIA0_9
timestamp 1681620392
transform 1 0 3043 0 1 2570
box -10 -3 10 3
use M3_M2  M3_M2_655
timestamp 1681620392
transform 1 0 132 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_787
timestamp 1681620392
transform 1 0 84 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_704
timestamp 1681620392
transform 1 0 84 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_856
timestamp 1681620392
transform 1 0 132 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_705
timestamp 1681620392
transform 1 0 156 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_745
timestamp 1681620392
transform 1 0 116 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_656
timestamp 1681620392
transform 1 0 204 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_788
timestamp 1681620392
transform 1 0 188 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_682
timestamp 1681620392
transform 1 0 196 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_789
timestamp 1681620392
transform 1 0 204 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_790
timestamp 1681620392
transform 1 0 220 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_683
timestamp 1681620392
transform 1 0 244 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_857
timestamp 1681620392
transform 1 0 188 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1681620392
transform 1 0 196 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1681620392
transform 1 0 212 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_860
timestamp 1681620392
transform 1 0 228 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_861
timestamp 1681620392
transform 1 0 236 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1681620392
transform 1 0 244 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_732
timestamp 1681620392
transform 1 0 196 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_746
timestamp 1681620392
transform 1 0 188 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_747
timestamp 1681620392
transform 1 0 212 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_863
timestamp 1681620392
transform 1 0 252 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_864
timestamp 1681620392
transform 1 0 260 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_748
timestamp 1681620392
transform 1 0 252 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_865
timestamp 1681620392
transform 1 0 284 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_657
timestamp 1681620392
transform 1 0 388 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_791
timestamp 1681620392
transform 1 0 388 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_866
timestamp 1681620392
transform 1 0 364 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_733
timestamp 1681620392
transform 1 0 364 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_867
timestamp 1681620392
transform 1 0 404 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_734
timestamp 1681620392
transform 1 0 404 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_658
timestamp 1681620392
transform 1 0 508 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_792
timestamp 1681620392
transform 1 0 508 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_868
timestamp 1681620392
transform 1 0 420 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_869
timestamp 1681620392
transform 1 0 476 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_684
timestamp 1681620392
transform 1 0 524 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_870
timestamp 1681620392
transform 1 0 524 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_749
timestamp 1681620392
transform 1 0 524 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_642
timestamp 1681620392
transform 1 0 620 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_659
timestamp 1681620392
transform 1 0 572 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_660
timestamp 1681620392
transform 1 0 612 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_793
timestamp 1681620392
transform 1 0 612 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_794
timestamp 1681620392
transform 1 0 628 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_871
timestamp 1681620392
transform 1 0 588 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_706
timestamp 1681620392
transform 1 0 612 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_643
timestamp 1681620392
transform 1 0 660 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_795
timestamp 1681620392
transform 1 0 652 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1681620392
transform 1 0 636 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_707
timestamp 1681620392
transform 1 0 652 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_796
timestamp 1681620392
transform 1 0 660 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_685
timestamp 1681620392
transform 1 0 668 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_708
timestamp 1681620392
transform 1 0 668 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_942
timestamp 1681620392
transform 1 0 660 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_943
timestamp 1681620392
transform 1 0 668 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_797
timestamp 1681620392
transform 1 0 700 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_686
timestamp 1681620392
transform 1 0 708 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_687
timestamp 1681620392
transform 1 0 732 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_798
timestamp 1681620392
transform 1 0 796 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_873
timestamp 1681620392
transform 1 0 708 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1681620392
transform 1 0 716 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_875
timestamp 1681620392
transform 1 0 772 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_735
timestamp 1681620392
transform 1 0 716 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_736
timestamp 1681620392
transform 1 0 748 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_876
timestamp 1681620392
transform 1 0 812 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_661
timestamp 1681620392
transform 1 0 844 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_662
timestamp 1681620392
transform 1 0 868 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_799
timestamp 1681620392
transform 1 0 844 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_877
timestamp 1681620392
transform 1 0 836 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_800
timestamp 1681620392
transform 1 0 964 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1681620392
transform 1 0 860 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_737
timestamp 1681620392
transform 1 0 844 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_944
timestamp 1681620392
transform 1 0 852 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_750
timestamp 1681620392
transform 1 0 836 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_960
timestamp 1681620392
transform 1 0 844 0 1 2505
box -2 -2 2 2
use M3_M2  M3_M2_751
timestamp 1681620392
transform 1 0 852 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_709
timestamp 1681620392
transform 1 0 876 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_879
timestamp 1681620392
transform 1 0 884 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_880
timestamp 1681620392
transform 1 0 940 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_945
timestamp 1681620392
transform 1 0 876 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_663
timestamp 1681620392
transform 1 0 980 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_801
timestamp 1681620392
transform 1 0 980 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_802
timestamp 1681620392
transform 1 0 996 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_881
timestamp 1681620392
transform 1 0 996 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_786
timestamp 1681620392
transform 1 0 1012 0 1 2545
box -2 -2 2 2
use M3_M2  M3_M2_688
timestamp 1681620392
transform 1 0 1012 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_803
timestamp 1681620392
transform 1 0 1020 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_710
timestamp 1681620392
transform 1 0 1052 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_882
timestamp 1681620392
transform 1 0 1060 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_883
timestamp 1681620392
transform 1 0 1076 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_752
timestamp 1681620392
transform 1 0 1076 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_644
timestamp 1681620392
transform 1 0 1092 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_689
timestamp 1681620392
transform 1 0 1092 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_884
timestamp 1681620392
transform 1 0 1092 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_711
timestamp 1681620392
transform 1 0 1100 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_885
timestamp 1681620392
transform 1 0 1132 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_738
timestamp 1681620392
transform 1 0 1132 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_664
timestamp 1681620392
transform 1 0 1156 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_804
timestamp 1681620392
transform 1 0 1156 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_805
timestamp 1681620392
transform 1 0 1164 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_753
timestamp 1681620392
transform 1 0 1164 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_665
timestamp 1681620392
transform 1 0 1204 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_806
timestamp 1681620392
transform 1 0 1204 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_886
timestamp 1681620392
transform 1 0 1180 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1681620392
transform 1 0 1196 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_739
timestamp 1681620392
transform 1 0 1180 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_690
timestamp 1681620392
transform 1 0 1220 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_807
timestamp 1681620392
transform 1 0 1228 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_712
timestamp 1681620392
transform 1 0 1212 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_888
timestamp 1681620392
transform 1 0 1228 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_889
timestamp 1681620392
transform 1 0 1244 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_946
timestamp 1681620392
transform 1 0 1228 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_691
timestamp 1681620392
transform 1 0 1268 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_645
timestamp 1681620392
transform 1 0 1356 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_666
timestamp 1681620392
transform 1 0 1324 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_808
timestamp 1681620392
transform 1 0 1356 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1681620392
transform 1 0 1268 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_891
timestamp 1681620392
transform 1 0 1276 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1681620392
transform 1 0 1332 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_740
timestamp 1681620392
transform 1 0 1316 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_741
timestamp 1681620392
transform 1 0 1332 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_667
timestamp 1681620392
transform 1 0 1380 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_809
timestamp 1681620392
transform 1 0 1380 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_947
timestamp 1681620392
transform 1 0 1404 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_810
timestamp 1681620392
transform 1 0 1428 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_713
timestamp 1681620392
transform 1 0 1428 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_893
timestamp 1681620392
transform 1 0 1444 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1681620392
transform 1 0 1436 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_811
timestamp 1681620392
transform 1 0 1484 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_812
timestamp 1681620392
transform 1 0 1492 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_813
timestamp 1681620392
transform 1 0 1516 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_714
timestamp 1681620392
transform 1 0 1484 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1681620392
transform 1 0 1508 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_716
timestamp 1681620392
transform 1 0 1524 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_742
timestamp 1681620392
transform 1 0 1516 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_814
timestamp 1681620392
transform 1 0 1540 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_717
timestamp 1681620392
transform 1 0 1540 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_668
timestamp 1681620392
transform 1 0 1572 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_669
timestamp 1681620392
transform 1 0 1612 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_815
timestamp 1681620392
transform 1 0 1572 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_816
timestamp 1681620392
transform 1 0 1588 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_894
timestamp 1681620392
transform 1 0 1556 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_692
timestamp 1681620392
transform 1 0 1620 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_631
timestamp 1681620392
transform 1 0 1700 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_817
timestamp 1681620392
transform 1 0 1684 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_818
timestamp 1681620392
transform 1 0 1692 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_895
timestamp 1681620392
transform 1 0 1612 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_718
timestamp 1681620392
transform 1 0 1660 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_632
timestamp 1681620392
transform 1 0 1764 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_633
timestamp 1681620392
transform 1 0 1836 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_634
timestamp 1681620392
transform 1 0 1852 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_635
timestamp 1681620392
transform 1 0 1868 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_670
timestamp 1681620392
transform 1 0 1748 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_671
timestamp 1681620392
transform 1 0 1788 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_819
timestamp 1681620392
transform 1 0 1716 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_820
timestamp 1681620392
transform 1 0 1724 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_821
timestamp 1681620392
transform 1 0 1748 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_822
timestamp 1681620392
transform 1 0 1764 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_896
timestamp 1681620392
transform 1 0 1668 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_897
timestamp 1681620392
transform 1 0 1676 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_898
timestamp 1681620392
transform 1 0 1692 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_899
timestamp 1681620392
transform 1 0 1700 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_900
timestamp 1681620392
transform 1 0 1716 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_949
timestamp 1681620392
transform 1 0 1572 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_754
timestamp 1681620392
transform 1 0 1556 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_755
timestamp 1681620392
transform 1 0 1580 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_743
timestamp 1681620392
transform 1 0 1684 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_756
timestamp 1681620392
transform 1 0 1692 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_770
timestamp 1681620392
transform 1 0 1668 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_719
timestamp 1681620392
transform 1 0 1724 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_950
timestamp 1681620392
transform 1 0 1716 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_744
timestamp 1681620392
transform 1 0 1724 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_693
timestamp 1681620392
transform 1 0 1844 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_823
timestamp 1681620392
transform 1 0 1852 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_636
timestamp 1681620392
transform 1 0 1932 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_646
timestamp 1681620392
transform 1 0 1908 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_672
timestamp 1681620392
transform 1 0 1892 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_673
timestamp 1681620392
transform 1 0 1916 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_824
timestamp 1681620392
transform 1 0 1876 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_694
timestamp 1681620392
transform 1 0 1884 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_825
timestamp 1681620392
transform 1 0 1892 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_826
timestamp 1681620392
transform 1 0 1900 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_901
timestamp 1681620392
transform 1 0 1788 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1681620392
transform 1 0 1844 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_903
timestamp 1681620392
transform 1 0 1852 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_951
timestamp 1681620392
transform 1 0 1748 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_720
timestamp 1681620392
transform 1 0 1868 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_904
timestamp 1681620392
transform 1 0 1876 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_757
timestamp 1681620392
transform 1 0 1812 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_758
timestamp 1681620392
transform 1 0 1852 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_952
timestamp 1681620392
transform 1 0 1876 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_721
timestamp 1681620392
transform 1 0 1892 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_827
timestamp 1681620392
transform 1 0 1924 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_905
timestamp 1681620392
transform 1 0 1908 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_722
timestamp 1681620392
transform 1 0 1924 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_647
timestamp 1681620392
transform 1 0 1948 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_674
timestamp 1681620392
transform 1 0 1940 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_828
timestamp 1681620392
transform 1 0 1940 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_829
timestamp 1681620392
transform 1 0 1948 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_906
timestamp 1681620392
transform 1 0 1932 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_953
timestamp 1681620392
transform 1 0 1924 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_675
timestamp 1681620392
transform 1 0 1988 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_695
timestamp 1681620392
transform 1 0 1956 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_830
timestamp 1681620392
transform 1 0 1964 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_696
timestamp 1681620392
transform 1 0 1980 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_831
timestamp 1681620392
transform 1 0 1988 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_697
timestamp 1681620392
transform 1 0 2004 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_907
timestamp 1681620392
transform 1 0 1956 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_908
timestamp 1681620392
transform 1 0 1964 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_909
timestamp 1681620392
transform 1 0 1980 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_910
timestamp 1681620392
transform 1 0 1996 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_911
timestamp 1681620392
transform 1 0 2004 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_759
timestamp 1681620392
transform 1 0 1956 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_760
timestamp 1681620392
transform 1 0 1996 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_776
timestamp 1681620392
transform 1 0 1980 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_832
timestamp 1681620392
transform 1 0 2020 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_833
timestamp 1681620392
transform 1 0 2052 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_912
timestamp 1681620392
transform 1 0 2036 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_723
timestamp 1681620392
transform 1 0 2044 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_913
timestamp 1681620392
transform 1 0 2052 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_761
timestamp 1681620392
transform 1 0 2052 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_771
timestamp 1681620392
transform 1 0 2020 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_772
timestamp 1681620392
transform 1 0 2036 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_834
timestamp 1681620392
transform 1 0 2068 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_835
timestamp 1681620392
transform 1 0 2084 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_914
timestamp 1681620392
transform 1 0 2076 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_773
timestamp 1681620392
transform 1 0 2076 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_698
timestamp 1681620392
transform 1 0 2108 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_637
timestamp 1681620392
transform 1 0 2148 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_638
timestamp 1681620392
transform 1 0 2172 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_639
timestamp 1681620392
transform 1 0 2244 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_640
timestamp 1681620392
transform 1 0 2260 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_676
timestamp 1681620392
transform 1 0 2140 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_836
timestamp 1681620392
transform 1 0 2116 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_837
timestamp 1681620392
transform 1 0 2148 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_915
timestamp 1681620392
transform 1 0 2100 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_916
timestamp 1681620392
transform 1 0 2108 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_917
timestamp 1681620392
transform 1 0 2124 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_918
timestamp 1681620392
transform 1 0 2140 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_954
timestamp 1681620392
transform 1 0 2100 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_774
timestamp 1681620392
transform 1 0 2100 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_762
timestamp 1681620392
transform 1 0 2140 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_648
timestamp 1681620392
transform 1 0 2244 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_838
timestamp 1681620392
transform 1 0 2244 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_839
timestamp 1681620392
transform 1 0 2260 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_919
timestamp 1681620392
transform 1 0 2156 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1681620392
transform 1 0 2164 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_921
timestamp 1681620392
transform 1 0 2204 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_724
timestamp 1681620392
transform 1 0 2244 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_763
timestamp 1681620392
transform 1 0 2156 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_764
timestamp 1681620392
transform 1 0 2180 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_765
timestamp 1681620392
transform 1 0 2212 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_641
timestamp 1681620392
transform 1 0 2364 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_649
timestamp 1681620392
transform 1 0 2292 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_840
timestamp 1681620392
transform 1 0 2292 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_841
timestamp 1681620392
transform 1 0 2380 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_922
timestamp 1681620392
transform 1 0 2276 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1681620392
transform 1 0 2324 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_725
timestamp 1681620392
transform 1 0 2356 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_650
timestamp 1681620392
transform 1 0 2420 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_842
timestamp 1681620392
transform 1 0 2420 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_699
timestamp 1681620392
transform 1 0 2460 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_700
timestamp 1681620392
transform 1 0 2492 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_651
timestamp 1681620392
transform 1 0 2516 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_843
timestamp 1681620392
transform 1 0 2516 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_701
timestamp 1681620392
transform 1 0 2588 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_924
timestamp 1681620392
transform 1 0 2372 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_925
timestamp 1681620392
transform 1 0 2388 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_926
timestamp 1681620392
transform 1 0 2404 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1681620392
transform 1 0 2444 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_928
timestamp 1681620392
transform 1 0 2500 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_955
timestamp 1681620392
transform 1 0 2276 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_766
timestamp 1681620392
transform 1 0 2316 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_767
timestamp 1681620392
transform 1 0 2372 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_775
timestamp 1681620392
transform 1 0 2276 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_777
timestamp 1681620392
transform 1 0 2388 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_778
timestamp 1681620392
transform 1 0 2476 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_726
timestamp 1681620392
transform 1 0 2516 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_929
timestamp 1681620392
transform 1 0 2540 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_727
timestamp 1681620392
transform 1 0 2548 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_652
timestamp 1681620392
transform 1 0 2612 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_930
timestamp 1681620392
transform 1 0 2596 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_956
timestamp 1681620392
transform 1 0 2604 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_677
timestamp 1681620392
transform 1 0 2628 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_844
timestamp 1681620392
transform 1 0 2620 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_931
timestamp 1681620392
transform 1 0 2620 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_932
timestamp 1681620392
transform 1 0 2636 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_957
timestamp 1681620392
transform 1 0 2628 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_845
timestamp 1681620392
transform 1 0 2652 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_933
timestamp 1681620392
transform 1 0 2660 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_846
timestamp 1681620392
transform 1 0 2684 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_702
timestamp 1681620392
transform 1 0 2692 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_678
timestamp 1681620392
transform 1 0 2724 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_847
timestamp 1681620392
transform 1 0 2716 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_848
timestamp 1681620392
transform 1 0 2724 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_934
timestamp 1681620392
transform 1 0 2692 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_935
timestamp 1681620392
transform 1 0 2708 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_728
timestamp 1681620392
transform 1 0 2716 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_653
timestamp 1681620392
transform 1 0 2748 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_654
timestamp 1681620392
transform 1 0 2764 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_679
timestamp 1681620392
transform 1 0 2788 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_849
timestamp 1681620392
transform 1 0 2748 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_850
timestamp 1681620392
transform 1 0 2764 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_851
timestamp 1681620392
transform 1 0 2852 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1681620392
transform 1 0 2868 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_936
timestamp 1681620392
transform 1 0 2740 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_958
timestamp 1681620392
transform 1 0 2716 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_937
timestamp 1681620392
transform 1 0 2788 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_729
timestamp 1681620392
transform 1 0 2836 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_938
timestamp 1681620392
transform 1 0 2844 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_939
timestamp 1681620392
transform 1 0 2852 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_768
timestamp 1681620392
transform 1 0 2748 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_769
timestamp 1681620392
transform 1 0 2852 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_680
timestamp 1681620392
transform 1 0 2900 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_681
timestamp 1681620392
transform 1 0 2956 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_853
timestamp 1681620392
transform 1 0 2900 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_854
timestamp 1681620392
transform 1 0 2916 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_855
timestamp 1681620392
transform 1 0 2932 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_703
timestamp 1681620392
transform 1 0 3012 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_730
timestamp 1681620392
transform 1 0 2916 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_940
timestamp 1681620392
transform 1 0 2956 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_731
timestamp 1681620392
transform 1 0 3004 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_941
timestamp 1681620392
transform 1 0 3012 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_959
timestamp 1681620392
transform 1 0 2900 0 1 2515
box -2 -2 2 2
use Project_Top_VIA0  Project_Top_VIA0_10
timestamp 1681620392
transform 1 0 24 0 1 2470
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_41
timestamp 1681620392
transform 1 0 72 0 -1 2570
box -8 -3 104 105
use INVX2  INVX2_37
timestamp 1681620392
transform 1 0 168 0 -1 2570
box -9 -3 26 105
use OAI22X1  OAI22X1_6
timestamp 1681620392
transform 1 0 184 0 -1 2570
box -8 -3 46 105
use INVX2  INVX2_39
timestamp 1681620392
transform -1 0 240 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_40
timestamp 1681620392
transform -1 0 256 0 -1 2570
box -9 -3 26 105
use FILL  FILL_140
timestamp 1681620392
transform 1 0 256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_141
timestamp 1681620392
transform 1 0 264 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_41
timestamp 1681620392
transform -1 0 288 0 -1 2570
box -9 -3 26 105
use FILL  FILL_142
timestamp 1681620392
transform 1 0 288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_143
timestamp 1681620392
transform 1 0 296 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_42
timestamp 1681620392
transform -1 0 400 0 -1 2570
box -8 -3 104 105
use FILL  FILL_144
timestamp 1681620392
transform 1 0 400 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_42
timestamp 1681620392
transform -1 0 424 0 -1 2570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_43
timestamp 1681620392
transform -1 0 520 0 -1 2570
box -8 -3 104 105
use FILL  FILL_145
timestamp 1681620392
transform 1 0 520 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_44
timestamp 1681620392
transform -1 0 624 0 -1 2570
box -8 -3 104 105
use OAI21X1  OAI21X1_45
timestamp 1681620392
transform 1 0 624 0 -1 2570
box -8 -3 34 105
use FILL  FILL_147
timestamp 1681620392
transform 1 0 656 0 -1 2570
box -8 -3 16 105
use FILL  FILL_151
timestamp 1681620392
transform 1 0 664 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_46
timestamp 1681620392
transform -1 0 704 0 -1 2570
box -8 -3 34 105
use FILL  FILL_152
timestamp 1681620392
transform 1 0 704 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1681620392
transform -1 0 808 0 -1 2570
box -8 -3 104 105
use FILL  FILL_155
timestamp 1681620392
transform 1 0 808 0 -1 2570
box -8 -3 16 105
use AND2X2  AND2X2_0
timestamp 1681620392
transform -1 0 848 0 -1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_18
timestamp 1681620392
transform 1 0 848 0 -1 2570
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_49
timestamp 1681620392
transform -1 0 976 0 -1 2570
box -8 -3 104 105
use FILL  FILL_156
timestamp 1681620392
transform 1 0 976 0 -1 2570
box -8 -3 16 105
use FILL  FILL_157
timestamp 1681620392
transform 1 0 984 0 -1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_12
timestamp 1681620392
transform -1 0 1016 0 -1 2570
box -8 -3 32 105
use OR2X1  OR2X1_1
timestamp 1681620392
transform 1 0 1016 0 -1 2570
box -8 -3 40 105
use INVX2  INVX2_44
timestamp 1681620392
transform 1 0 1048 0 -1 2570
box -9 -3 26 105
use FILL  FILL_158
timestamp 1681620392
transform 1 0 1064 0 -1 2570
box -8 -3 16 105
use FILL  FILL_159
timestamp 1681620392
transform 1 0 1072 0 -1 2570
box -8 -3 16 105
use FILL  FILL_160
timestamp 1681620392
transform 1 0 1080 0 -1 2570
box -8 -3 16 105
use FILL  FILL_161
timestamp 1681620392
transform 1 0 1088 0 -1 2570
box -8 -3 16 105
use FILL  FILL_162
timestamp 1681620392
transform 1 0 1096 0 -1 2570
box -8 -3 16 105
use FILL  FILL_163
timestamp 1681620392
transform 1 0 1104 0 -1 2570
box -8 -3 16 105
use AND2X2  AND2X2_1
timestamp 1681620392
transform -1 0 1144 0 -1 2570
box -8 -3 40 105
use FILL  FILL_165
timestamp 1681620392
transform 1 0 1144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_166
timestamp 1681620392
transform 1 0 1152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_167
timestamp 1681620392
transform 1 0 1160 0 -1 2570
box -8 -3 16 105
use AND2X2  AND2X2_2
timestamp 1681620392
transform 1 0 1168 0 -1 2570
box -8 -3 40 105
use FILL  FILL_168
timestamp 1681620392
transform 1 0 1200 0 -1 2570
box -8 -3 16 105
use NAND2X1  NAND2X1_29
timestamp 1681620392
transform 1 0 1208 0 -1 2570
box -8 -3 32 105
use AND2X2  AND2X2_3
timestamp 1681620392
transform 1 0 1232 0 -1 2570
box -8 -3 40 105
use FILL  FILL_174
timestamp 1681620392
transform 1 0 1264 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_50
timestamp 1681620392
transform -1 0 1368 0 -1 2570
box -8 -3 104 105
use FILL  FILL_175
timestamp 1681620392
transform 1 0 1368 0 -1 2570
box -8 -3 16 105
use FILL  FILL_176
timestamp 1681620392
transform 1 0 1376 0 -1 2570
box -8 -3 16 105
use FILL  FILL_177
timestamp 1681620392
transform 1 0 1384 0 -1 2570
box -8 -3 16 105
use FILL  FILL_178
timestamp 1681620392
transform 1 0 1392 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_53
timestamp 1681620392
transform -1 0 1432 0 -1 2570
box -8 -3 34 105
use FILL  FILL_179
timestamp 1681620392
transform 1 0 1432 0 -1 2570
box -8 -3 16 105
use FILL  FILL_180
timestamp 1681620392
transform 1 0 1440 0 -1 2570
box -8 -3 16 105
use FILL  FILL_182
timestamp 1681620392
transform 1 0 1448 0 -1 2570
box -8 -3 16 105
use FILL  FILL_187
timestamp 1681620392
transform 1 0 1456 0 -1 2570
box -8 -3 16 105
use NAND2X1  NAND2X1_34
timestamp 1681620392
transform -1 0 1488 0 -1 2570
box -8 -3 32 105
use OAI21X1  OAI21X1_56
timestamp 1681620392
transform -1 0 1520 0 -1 2570
box -8 -3 34 105
use FILL  FILL_188
timestamp 1681620392
transform 1 0 1520 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_47
timestamp 1681620392
transform -1 0 1544 0 -1 2570
box -9 -3 26 105
use M3_M2  M3_M2_779
timestamp 1681620392
transform 1 0 1556 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_780
timestamp 1681620392
transform 1 0 1572 0 1 2475
box -3 -3 3 3
use OAI21X1  OAI21X1_57
timestamp 1681620392
transform 1 0 1544 0 -1 2570
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_52
timestamp 1681620392
transform 1 0 1576 0 -1 2570
box -8 -3 104 105
use INVX2  INVX2_59
timestamp 1681620392
transform -1 0 1688 0 -1 2570
box -9 -3 26 105
use M3_M2  M3_M2_781
timestamp 1681620392
transform 1 0 1724 0 1 2475
box -3 -3 3 3
use OAI21X1  OAI21X1_67
timestamp 1681620392
transform 1 0 1688 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_68
timestamp 1681620392
transform 1 0 1720 0 -1 2570
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_57
timestamp 1681620392
transform 1 0 1752 0 -1 2570
box -8 -3 104 105
use OAI21X1  OAI21X1_69
timestamp 1681620392
transform 1 0 1848 0 -1 2570
box -8 -3 34 105
use INVX2  INVX2_60
timestamp 1681620392
transform -1 0 1896 0 -1 2570
box -9 -3 26 105
use OAI21X1  OAI21X1_70
timestamp 1681620392
transform 1 0 1896 0 -1 2570
box -8 -3 34 105
use INVX2  INVX2_61
timestamp 1681620392
transform -1 0 1944 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_62
timestamp 1681620392
transform 1 0 1944 0 -1 2570
box -9 -3 26 105
use AOI22X1  AOI22X1_15
timestamp 1681620392
transform 1 0 1960 0 -1 2570
box -8 -3 46 105
use FILL  FILL_205
timestamp 1681620392
transform 1 0 2000 0 -1 2570
box -8 -3 16 105
use FILL  FILL_206
timestamp 1681620392
transform 1 0 2008 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_16
timestamp 1681620392
transform 1 0 2016 0 -1 2570
box -8 -3 46 105
use INVX2  INVX2_63
timestamp 1681620392
transform -1 0 2072 0 -1 2570
box -9 -3 26 105
use FILL  FILL_207
timestamp 1681620392
transform 1 0 2072 0 -1 2570
box -8 -3 16 105
use NAND2X1  NAND2X1_37
timestamp 1681620392
transform 1 0 2080 0 -1 2570
box -8 -3 32 105
use M3_M2  M3_M2_782
timestamp 1681620392
transform 1 0 2116 0 1 2475
box -3 -3 3 3
use AOI22X1  AOI22X1_17
timestamp 1681620392
transform 1 0 2104 0 -1 2570
box -8 -3 46 105
use INVX2  INVX2_64
timestamp 1681620392
transform 1 0 2144 0 -1 2570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_58
timestamp 1681620392
transform -1 0 2256 0 -1 2570
box -8 -3 104 105
use NAND2X1  NAND2X1_38
timestamp 1681620392
transform 1 0 2256 0 -1 2570
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_59
timestamp 1681620392
transform 1 0 2280 0 -1 2570
box -8 -3 104 105
use AND2X2  AND2X2_4
timestamp 1681620392
transform 1 0 2376 0 -1 2570
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_60
timestamp 1681620392
transform 1 0 2408 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_61
timestamp 1681620392
transform 1 0 2504 0 -1 2570
box -8 -3 104 105
use NAND2X1  NAND2X1_39
timestamp 1681620392
transform -1 0 2624 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_40
timestamp 1681620392
transform -1 0 2648 0 -1 2570
box -8 -3 32 105
use FILL  FILL_208
timestamp 1681620392
transform 1 0 2648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_209
timestamp 1681620392
transform 1 0 2656 0 -1 2570
box -8 -3 16 105
use FILL  FILL_210
timestamp 1681620392
transform 1 0 2664 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_18
timestamp 1681620392
transform 1 0 2672 0 -1 2570
box -8 -3 46 105
use FILL  FILL_211
timestamp 1681620392
transform 1 0 2712 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_71
timestamp 1681620392
transform -1 0 2752 0 -1 2570
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_62
timestamp 1681620392
transform 1 0 2752 0 -1 2570
box -8 -3 104 105
use INVX2  INVX2_65
timestamp 1681620392
transform 1 0 2848 0 -1 2570
box -9 -3 26 105
use OAI21X1  OAI21X1_72
timestamp 1681620392
transform 1 0 2864 0 -1 2570
box -8 -3 34 105
use NAND2X1  NAND2X1_41
timestamp 1681620392
transform -1 0 2920 0 -1 2570
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_63
timestamp 1681620392
transform 1 0 2920 0 -1 2570
box -8 -3 104 105
use Project_Top_VIA0  Project_Top_VIA0_11
timestamp 1681620392
transform 1 0 3067 0 1 2470
box -10 -3 10 3
use M2_M1  M2_M1_1004
timestamp 1681620392
transform 1 0 132 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1076
timestamp 1681620392
transform 1 0 68 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_872
timestamp 1681620392
transform 1 0 132 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_808
timestamp 1681620392
transform 1 0 220 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_793
timestamp 1681620392
transform 1 0 252 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_961
timestamp 1681620392
transform 1 0 252 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_966
timestamp 1681620392
transform 1 0 196 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_967
timestamp 1681620392
transform 1 0 204 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_968
timestamp 1681620392
transform 1 0 236 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1005
timestamp 1681620392
transform 1 0 180 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1077
timestamp 1681620392
transform 1 0 156 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1078
timestamp 1681620392
transform 1 0 172 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_873
timestamp 1681620392
transform 1 0 188 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_1006
timestamp 1681620392
transform 1 0 220 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1079
timestamp 1681620392
transform 1 0 196 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_891
timestamp 1681620392
transform 1 0 196 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_892
timestamp 1681620392
transform 1 0 212 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_794
timestamp 1681620392
transform 1 0 276 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_809
timestamp 1681620392
transform 1 0 284 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_969
timestamp 1681620392
transform 1 0 260 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_854
timestamp 1681620392
transform 1 0 260 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_970
timestamp 1681620392
transform 1 0 292 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_810
timestamp 1681620392
transform 1 0 324 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_832
timestamp 1681620392
transform 1 0 316 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_1007
timestamp 1681620392
transform 1 0 284 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1080
timestamp 1681620392
transform 1 0 244 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_855
timestamp 1681620392
transform 1 0 292 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_856
timestamp 1681620392
transform 1 0 308 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_1008
timestamp 1681620392
transform 1 0 316 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1009
timestamp 1681620392
transform 1 0 324 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_874
timestamp 1681620392
transform 1 0 276 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_1081
timestamp 1681620392
transform 1 0 284 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1082
timestamp 1681620392
transform 1 0 292 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_893
timestamp 1681620392
transform 1 0 244 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_894
timestamp 1681620392
transform 1 0 260 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_1152
timestamp 1681620392
transform 1 0 268 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_895
timestamp 1681620392
transform 1 0 284 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_833
timestamp 1681620392
transform 1 0 340 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_811
timestamp 1681620392
transform 1 0 380 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_971
timestamp 1681620392
transform 1 0 364 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1010
timestamp 1681620392
transform 1 0 340 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_857
timestamp 1681620392
transform 1 0 356 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_1011
timestamp 1681620392
transform 1 0 364 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1083
timestamp 1681620392
transform 1 0 316 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1084
timestamp 1681620392
transform 1 0 332 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_875
timestamp 1681620392
transform 1 0 340 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_1085
timestamp 1681620392
transform 1 0 348 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1153
timestamp 1681620392
transform 1 0 340 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_896
timestamp 1681620392
transform 1 0 348 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_925
timestamp 1681620392
transform 1 0 332 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_876
timestamp 1681620392
transform 1 0 372 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_1086
timestamp 1681620392
transform 1 0 380 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_897
timestamp 1681620392
transform 1 0 388 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_1012
timestamp 1681620392
transform 1 0 404 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1087
timestamp 1681620392
transform 1 0 404 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_877
timestamp 1681620392
transform 1 0 412 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_1154
timestamp 1681620392
transform 1 0 412 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1088
timestamp 1681620392
transform 1 0 428 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_962
timestamp 1681620392
transform 1 0 444 0 1 2435
box -2 -2 2 2
use M3_M2  M3_M2_812
timestamp 1681620392
transform 1 0 452 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_972
timestamp 1681620392
transform 1 0 452 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1013
timestamp 1681620392
transform 1 0 452 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_878
timestamp 1681620392
transform 1 0 452 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_926
timestamp 1681620392
transform 1 0 444 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_927
timestamp 1681620392
transform 1 0 468 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_795
timestamp 1681620392
transform 1 0 572 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_813
timestamp 1681620392
transform 1 0 492 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_814
timestamp 1681620392
transform 1 0 532 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_973
timestamp 1681620392
transform 1 0 484 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_834
timestamp 1681620392
transform 1 0 548 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_1014
timestamp 1681620392
transform 1 0 492 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1015
timestamp 1681620392
transform 1 0 548 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1089
timestamp 1681620392
transform 1 0 572 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_835
timestamp 1681620392
transform 1 0 588 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_1016
timestamp 1681620392
transform 1 0 588 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_815
timestamp 1681620392
transform 1 0 604 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_1017
timestamp 1681620392
transform 1 0 604 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1090
timestamp 1681620392
transform 1 0 612 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_816
timestamp 1681620392
transform 1 0 716 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_963
timestamp 1681620392
transform 1 0 724 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_1018
timestamp 1681620392
transform 1 0 684 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_858
timestamp 1681620392
transform 1 0 708 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_1091
timestamp 1681620392
transform 1 0 708 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_898
timestamp 1681620392
transform 1 0 684 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_928
timestamp 1681620392
transform 1 0 644 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_929
timestamp 1681620392
transform 1 0 708 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_817
timestamp 1681620392
transform 1 0 732 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_974
timestamp 1681620392
transform 1 0 724 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1681620392
transform 1 0 732 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_836
timestamp 1681620392
transform 1 0 740 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_1019
timestamp 1681620392
transform 1 0 740 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_837
timestamp 1681620392
transform 1 0 788 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_1020
timestamp 1681620392
transform 1 0 780 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1021
timestamp 1681620392
transform 1 0 788 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1092
timestamp 1681620392
transform 1 0 764 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_879
timestamp 1681620392
transform 1 0 772 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_859
timestamp 1681620392
transform 1 0 796 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_1093
timestamp 1681620392
transform 1 0 788 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_899
timestamp 1681620392
transform 1 0 764 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_1094
timestamp 1681620392
transform 1 0 820 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_818
timestamp 1681620392
transform 1 0 836 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_964
timestamp 1681620392
transform 1 0 860 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_976
timestamp 1681620392
transform 1 0 836 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_977
timestamp 1681620392
transform 1 0 868 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_978
timestamp 1681620392
transform 1 0 876 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1022
timestamp 1681620392
transform 1 0 852 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_860
timestamp 1681620392
transform 1 0 868 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_965
timestamp 1681620392
transform 1 0 924 0 1 2435
box -2 -2 2 2
use M3_M2  M3_M2_838
timestamp 1681620392
transform 1 0 900 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_979
timestamp 1681620392
transform 1 0 908 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_839
timestamp 1681620392
transform 1 0 924 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_1023
timestamp 1681620392
transform 1 0 892 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_880
timestamp 1681620392
transform 1 0 868 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_1095
timestamp 1681620392
transform 1 0 876 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_861
timestamp 1681620392
transform 1 0 900 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_1024
timestamp 1681620392
transform 1 0 916 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1096
timestamp 1681620392
transform 1 0 900 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_930
timestamp 1681620392
transform 1 0 892 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_980
timestamp 1681620392
transform 1 0 940 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1097
timestamp 1681620392
transform 1 0 940 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_783
timestamp 1681620392
transform 1 0 964 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_900
timestamp 1681620392
transform 1 0 956 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_1025
timestamp 1681620392
transform 1 0 988 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1026
timestamp 1681620392
transform 1 0 996 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1098
timestamp 1681620392
transform 1 0 980 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_881
timestamp 1681620392
transform 1 0 988 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_901
timestamp 1681620392
transform 1 0 980 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_1099
timestamp 1681620392
transform 1 0 1012 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_840
timestamp 1681620392
transform 1 0 1028 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_1027
timestamp 1681620392
transform 1 0 1028 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_882
timestamp 1681620392
transform 1 0 1028 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_1100
timestamp 1681620392
transform 1 0 1052 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1155
timestamp 1681620392
transform 1 0 1028 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1156
timestamp 1681620392
transform 1 0 1036 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1028
timestamp 1681620392
transform 1 0 1076 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1029
timestamp 1681620392
transform 1 0 1148 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1101
timestamp 1681620392
transform 1 0 1100 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_902
timestamp 1681620392
transform 1 0 1148 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_819
timestamp 1681620392
transform 1 0 1212 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_981
timestamp 1681620392
transform 1 0 1212 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1030
timestamp 1681620392
transform 1 0 1212 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1031
timestamp 1681620392
transform 1 0 1228 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1102
timestamp 1681620392
transform 1 0 1212 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_903
timestamp 1681620392
transform 1 0 1212 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_1103
timestamp 1681620392
transform 1 0 1236 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1157
timestamp 1681620392
transform 1 0 1244 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_820
timestamp 1681620392
transform 1 0 1268 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_1032
timestamp 1681620392
transform 1 0 1276 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1104
timestamp 1681620392
transform 1 0 1284 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_931
timestamp 1681620392
transform 1 0 1260 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_796
timestamp 1681620392
transform 1 0 1308 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_1033
timestamp 1681620392
transform 1 0 1300 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_932
timestamp 1681620392
transform 1 0 1300 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_787
timestamp 1681620392
transform 1 0 1356 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_841
timestamp 1681620392
transform 1 0 1332 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_1034
timestamp 1681620392
transform 1 0 1332 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1035
timestamp 1681620392
transform 1 0 1380 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1036
timestamp 1681620392
transform 1 0 1428 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1105
timestamp 1681620392
transform 1 0 1324 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1158
timestamp 1681620392
transform 1 0 1316 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1681620392
transform 1 0 1348 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_904
timestamp 1681620392
transform 1 0 1348 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_905
timestamp 1681620392
transform 1 0 1396 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_906
timestamp 1681620392
transform 1 0 1420 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_862
timestamp 1681620392
transform 1 0 1444 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_821
timestamp 1681620392
transform 1 0 1548 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_842
timestamp 1681620392
transform 1 0 1540 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_982
timestamp 1681620392
transform 1 0 1548 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1037
timestamp 1681620392
transform 1 0 1492 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1038
timestamp 1681620392
transform 1 0 1524 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1107
timestamp 1681620392
transform 1 0 1444 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1108
timestamp 1681620392
transform 1 0 1532 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_907
timestamp 1681620392
transform 1 0 1444 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_797
timestamp 1681620392
transform 1 0 1572 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_798
timestamp 1681620392
transform 1 0 1596 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_983
timestamp 1681620392
transform 1 0 1572 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_843
timestamp 1681620392
transform 1 0 1588 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_1039
timestamp 1681620392
transform 1 0 1556 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1040
timestamp 1681620392
transform 1 0 1564 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1109
timestamp 1681620392
transform 1 0 1548 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_863
timestamp 1681620392
transform 1 0 1572 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_1041
timestamp 1681620392
transform 1 0 1580 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1110
timestamp 1681620392
transform 1 0 1572 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_933
timestamp 1681620392
transform 1 0 1564 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_822
timestamp 1681620392
transform 1 0 1628 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_799
timestamp 1681620392
transform 1 0 1732 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_984
timestamp 1681620392
transform 1 0 1628 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1111
timestamp 1681620392
transform 1 0 1604 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1112
timestamp 1681620392
transform 1 0 1612 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_908
timestamp 1681620392
transform 1 0 1604 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_844
timestamp 1681620392
transform 1 0 1644 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_845
timestamp 1681620392
transform 1 0 1716 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_788
timestamp 1681620392
transform 1 0 1756 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_985
timestamp 1681620392
transform 1 0 1732 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1042
timestamp 1681620392
transform 1 0 1668 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_864
timestamp 1681620392
transform 1 0 1676 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_865
timestamp 1681620392
transform 1 0 1708 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_846
timestamp 1681620392
transform 1 0 1740 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_1043
timestamp 1681620392
transform 1 0 1724 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1044
timestamp 1681620392
transform 1 0 1740 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1113
timestamp 1681620392
transform 1 0 1644 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_909
timestamp 1681620392
transform 1 0 1668 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_866
timestamp 1681620392
transform 1 0 1748 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_1045
timestamp 1681620392
transform 1 0 1772 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1114
timestamp 1681620392
transform 1 0 1748 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1115
timestamp 1681620392
transform 1 0 1756 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_867
timestamp 1681620392
transform 1 0 1788 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_800
timestamp 1681620392
transform 1 0 1812 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_823
timestamp 1681620392
transform 1 0 1828 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_847
timestamp 1681620392
transform 1 0 1812 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_986
timestamp 1681620392
transform 1 0 1820 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_987
timestamp 1681620392
transform 1 0 1828 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1046
timestamp 1681620392
transform 1 0 1796 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1047
timestamp 1681620392
transform 1 0 1804 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1116
timestamp 1681620392
transform 1 0 1780 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1117
timestamp 1681620392
transform 1 0 1804 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_801
timestamp 1681620392
transform 1 0 1852 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_784
timestamp 1681620392
transform 1 0 1884 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_824
timestamp 1681620392
transform 1 0 1844 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_825
timestamp 1681620392
transform 1 0 1868 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_988
timestamp 1681620392
transform 1 0 1852 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_989
timestamp 1681620392
transform 1 0 1868 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1048
timestamp 1681620392
transform 1 0 1844 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_802
timestamp 1681620392
transform 1 0 1900 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_803
timestamp 1681620392
transform 1 0 1932 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_1049
timestamp 1681620392
transform 1 0 1876 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1681620392
transform 1 0 1892 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1681620392
transform 1 0 1852 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1119
timestamp 1681620392
transform 1 0 1868 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1120
timestamp 1681620392
transform 1 0 1876 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_883
timestamp 1681620392
transform 1 0 1892 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_826
timestamp 1681620392
transform 1 0 2020 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_990
timestamp 1681620392
transform 1 0 2020 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1051
timestamp 1681620392
transform 1 0 1940 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1052
timestamp 1681620392
transform 1 0 1996 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1053
timestamp 1681620392
transform 1 0 2012 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1121
timestamp 1681620392
transform 1 0 1900 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1122
timestamp 1681620392
transform 1 0 1916 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1123
timestamp 1681620392
transform 1 0 2004 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_910
timestamp 1681620392
transform 1 0 1876 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_911
timestamp 1681620392
transform 1 0 1940 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1681620392
transform 1 0 1916 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_1124
timestamp 1681620392
transform 1 0 2028 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_785
timestamp 1681620392
transform 1 0 2044 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_789
timestamp 1681620392
transform 1 0 2044 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_991
timestamp 1681620392
transform 1 0 2044 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_790
timestamp 1681620392
transform 1 0 2100 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_791
timestamp 1681620392
transform 1 0 2124 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_992
timestamp 1681620392
transform 1 0 2076 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1054
timestamp 1681620392
transform 1 0 2052 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1055
timestamp 1681620392
transform 1 0 2060 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1125
timestamp 1681620392
transform 1 0 2044 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_884
timestamp 1681620392
transform 1 0 2060 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_1056
timestamp 1681620392
transform 1 0 2084 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1057
timestamp 1681620392
transform 1 0 2116 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1058
timestamp 1681620392
transform 1 0 2188 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1126
timestamp 1681620392
transform 1 0 2076 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1127
timestamp 1681620392
transform 1 0 2164 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1128
timestamp 1681620392
transform 1 0 2180 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_912
timestamp 1681620392
transform 1 0 2076 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_913
timestamp 1681620392
transform 1 0 2116 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_914
timestamp 1681620392
transform 1 0 2164 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_885
timestamp 1681620392
transform 1 0 2188 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_804
timestamp 1681620392
transform 1 0 2268 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_827
timestamp 1681620392
transform 1 0 2228 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_828
timestamp 1681620392
transform 1 0 2252 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_993
timestamp 1681620392
transform 1 0 2228 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_994
timestamp 1681620392
transform 1 0 2252 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1059
timestamp 1681620392
transform 1 0 2244 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1060
timestamp 1681620392
transform 1 0 2252 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1129
timestamp 1681620392
transform 1 0 2204 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1130
timestamp 1681620392
transform 1 0 2212 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1131
timestamp 1681620392
transform 1 0 2228 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_935
timestamp 1681620392
transform 1 0 2172 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_886
timestamp 1681620392
transform 1 0 2252 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_936
timestamp 1681620392
transform 1 0 2228 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_1132
timestamp 1681620392
transform 1 0 2276 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1133
timestamp 1681620392
transform 1 0 2284 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_829
timestamp 1681620392
transform 1 0 2316 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_995
timestamp 1681620392
transform 1 0 2316 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_868
timestamp 1681620392
transform 1 0 2316 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_1134
timestamp 1681620392
transform 1 0 2324 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_848
timestamp 1681620392
transform 1 0 2364 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_1061
timestamp 1681620392
transform 1 0 2364 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1135
timestamp 1681620392
transform 1 0 2372 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1136
timestamp 1681620392
transform 1 0 2388 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_996
timestamp 1681620392
transform 1 0 2404 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_869
timestamp 1681620392
transform 1 0 2404 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_805
timestamp 1681620392
transform 1 0 2420 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_830
timestamp 1681620392
transform 1 0 2428 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_806
timestamp 1681620392
transform 1 0 2452 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_831
timestamp 1681620392
transform 1 0 2468 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_849
timestamp 1681620392
transform 1 0 2452 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_997
timestamp 1681620392
transform 1 0 2468 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1062
timestamp 1681620392
transform 1 0 2452 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1137
timestamp 1681620392
transform 1 0 2436 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1138
timestamp 1681620392
transform 1 0 2460 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_915
timestamp 1681620392
transform 1 0 2460 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_807
timestamp 1681620392
transform 1 0 2492 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_887
timestamp 1681620392
transform 1 0 2484 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_998
timestamp 1681620392
transform 1 0 2500 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1063
timestamp 1681620392
transform 1 0 2516 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1139
timestamp 1681620392
transform 1 0 2524 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_850
timestamp 1681620392
transform 1 0 2548 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_1064
timestamp 1681620392
transform 1 0 2548 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1140
timestamp 1681620392
transform 1 0 2532 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_792
timestamp 1681620392
transform 1 0 2564 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_999
timestamp 1681620392
transform 1 0 2564 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1065
timestamp 1681620392
transform 1 0 2564 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_916
timestamp 1681620392
transform 1 0 2556 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_1141
timestamp 1681620392
transform 1 0 2572 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_917
timestamp 1681620392
transform 1 0 2572 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_1066
timestamp 1681620392
transform 1 0 2604 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1681620392
transform 1 0 2588 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1143
timestamp 1681620392
transform 1 0 2596 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_918
timestamp 1681620392
transform 1 0 2604 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_937
timestamp 1681620392
transform 1 0 2596 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_870
timestamp 1681620392
transform 1 0 2644 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_786
timestamp 1681620392
transform 1 0 2668 0 1 2465
box -3 -3 3 3
use M2_M1  M2_M1_1000
timestamp 1681620392
transform 1 0 2676 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1681620392
transform 1 0 2652 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1068
timestamp 1681620392
transform 1 0 2668 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_888
timestamp 1681620392
transform 1 0 2636 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_889
timestamp 1681620392
transform 1 0 2652 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_871
timestamp 1681620392
transform 1 0 2676 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_1069
timestamp 1681620392
transform 1 0 2692 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1144
timestamp 1681620392
transform 1 0 2708 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_851
timestamp 1681620392
transform 1 0 2740 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_1070
timestamp 1681620392
transform 1 0 2732 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1071
timestamp 1681620392
transform 1 0 2740 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_890
timestamp 1681620392
transform 1 0 2732 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_1145
timestamp 1681620392
transform 1 0 2740 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1681620392
transform 1 0 2748 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_938
timestamp 1681620392
transform 1 0 2724 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_1072
timestamp 1681620392
transform 1 0 2780 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_919
timestamp 1681620392
transform 1 0 2780 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_1147
timestamp 1681620392
transform 1 0 2804 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_920
timestamp 1681620392
transform 1 0 2804 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_1001
timestamp 1681620392
transform 1 0 2836 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1002
timestamp 1681620392
transform 1 0 2852 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1681620392
transform 1 0 2828 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1073
timestamp 1681620392
transform 1 0 2876 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_921
timestamp 1681620392
transform 1 0 2868 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_1149
timestamp 1681620392
transform 1 0 2884 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1003
timestamp 1681620392
transform 1 0 2900 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_922
timestamp 1681620392
transform 1 0 2892 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_852
timestamp 1681620392
transform 1 0 2916 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_853
timestamp 1681620392
transform 1 0 3012 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_1074
timestamp 1681620392
transform 1 0 2956 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1075
timestamp 1681620392
transform 1 0 3012 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1150
timestamp 1681620392
transform 1 0 2916 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1151
timestamp 1681620392
transform 1 0 2932 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_923
timestamp 1681620392
transform 1 0 2916 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_924
timestamp 1681620392
transform 1 0 2956 0 1 2395
box -3 -3 3 3
use Project_Top_VIA0  Project_Top_VIA0_12
timestamp 1681620392
transform 1 0 48 0 1 2370
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_64
timestamp 1681620392
transform -1 0 168 0 1 2370
box -8 -3 104 105
use OAI21X1  OAI21X1_73
timestamp 1681620392
transform 1 0 168 0 1 2370
box -8 -3 34 105
use M3_M2  M3_M2_939
timestamp 1681620392
transform 1 0 236 0 1 2375
box -3 -3 3 3
use NAND3X1  NAND3X1_19
timestamp 1681620392
transform -1 0 232 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_20
timestamp 1681620392
transform 1 0 232 0 1 2370
box -8 -3 40 105
use NOR2X1  NOR2X1_15
timestamp 1681620392
transform 1 0 264 0 1 2370
box -8 -3 32 105
use OAI21X1  OAI21X1_74
timestamp 1681620392
transform -1 0 320 0 1 2370
box -8 -3 34 105
use NOR2X1  NOR2X1_16
timestamp 1681620392
transform -1 0 344 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_42
timestamp 1681620392
transform 1 0 344 0 1 2370
box -8 -3 32 105
use INVX2  INVX2_66
timestamp 1681620392
transform -1 0 384 0 1 2370
box -9 -3 26 105
use M3_M2  M3_M2_940
timestamp 1681620392
transform 1 0 404 0 1 2375
box -3 -3 3 3
use NOR2X1  NOR2X1_17
timestamp 1681620392
transform 1 0 384 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_18
timestamp 1681620392
transform 1 0 408 0 1 2370
box -8 -3 32 105
use FILL  FILL_212
timestamp 1681620392
transform 1 0 432 0 1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_21
timestamp 1681620392
transform 1 0 440 0 1 2370
box -8 -3 40 105
use FILL  FILL_213
timestamp 1681620392
transform 1 0 472 0 1 2370
box -8 -3 16 105
use FILL  FILL_221
timestamp 1681620392
transform 1 0 480 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_65
timestamp 1681620392
transform -1 0 584 0 1 2370
box -8 -3 104 105
use FILL  FILL_222
timestamp 1681620392
transform 1 0 584 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_71
timestamp 1681620392
transform -1 0 608 0 1 2370
box -9 -3 26 105
use FILL  FILL_223
timestamp 1681620392
transform 1 0 608 0 1 2370
box -8 -3 16 105
use FILL  FILL_224
timestamp 1681620392
transform 1 0 616 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_66
timestamp 1681620392
transform -1 0 720 0 1 2370
box -8 -3 104 105
use FILL  FILL_225
timestamp 1681620392
transform 1 0 720 0 1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_26
timestamp 1681620392
transform 1 0 728 0 1 2370
box -8 -3 40 105
use OAI21X1  OAI21X1_76
timestamp 1681620392
transform -1 0 792 0 1 2370
box -8 -3 34 105
use FILL  FILL_226
timestamp 1681620392
transform 1 0 792 0 1 2370
box -8 -3 16 105
use FILL  FILL_227
timestamp 1681620392
transform 1 0 800 0 1 2370
box -8 -3 16 105
use FILL  FILL_228
timestamp 1681620392
transform 1 0 808 0 1 2370
box -8 -3 16 105
use NAND2X1  NAND2X1_47
timestamp 1681620392
transform 1 0 816 0 1 2370
box -8 -3 32 105
use NAND3X1  NAND3X1_28
timestamp 1681620392
transform 1 0 840 0 1 2370
box -8 -3 40 105
use OAI21X1  OAI21X1_78
timestamp 1681620392
transform -1 0 904 0 1 2370
box -8 -3 34 105
use NAND3X1  NAND3X1_29
timestamp 1681620392
transform 1 0 904 0 1 2370
box -8 -3 40 105
use FILL  FILL_234
timestamp 1681620392
transform 1 0 936 0 1 2370
box -8 -3 16 105
use FILL  FILL_235
timestamp 1681620392
transform 1 0 944 0 1 2370
box -8 -3 16 105
use FILL  FILL_236
timestamp 1681620392
transform 1 0 952 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_73
timestamp 1681620392
transform 1 0 960 0 1 2370
box -9 -3 26 105
use FILL  FILL_237
timestamp 1681620392
transform 1 0 976 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_74
timestamp 1681620392
transform 1 0 984 0 1 2370
box -9 -3 26 105
use FILL  FILL_238
timestamp 1681620392
transform 1 0 1000 0 1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_20
timestamp 1681620392
transform -1 0 1032 0 1 2370
box -8 -3 32 105
use AOI21X1  AOI21X1_7
timestamp 1681620392
transform -1 0 1064 0 1 2370
box -7 -3 39 105
use FILL  FILL_239
timestamp 1681620392
transform 1 0 1064 0 1 2370
box -8 -3 16 105
use FILL  FILL_240
timestamp 1681620392
transform 1 0 1072 0 1 2370
box -8 -3 16 105
use FILL  FILL_241
timestamp 1681620392
transform 1 0 1080 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_941
timestamp 1681620392
transform 1 0 1180 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_69
timestamp 1681620392
transform 1 0 1088 0 1 2370
box -8 -3 104 105
use FILL  FILL_242
timestamp 1681620392
transform 1 0 1184 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_75
timestamp 1681620392
transform 1 0 1192 0 1 2370
box -9 -3 26 105
use M3_M2  M3_M2_942
timestamp 1681620392
transform 1 0 1244 0 1 2375
box -3 -3 3 3
use OAI21X1  OAI21X1_79
timestamp 1681620392
transform -1 0 1240 0 1 2370
box -8 -3 34 105
use FILL  FILL_243
timestamp 1681620392
transform 1 0 1240 0 1 2370
box -8 -3 16 105
use OR2X1  OR2X1_3
timestamp 1681620392
transform 1 0 1248 0 1 2370
box -8 -3 40 105
use M3_M2  M3_M2_943
timestamp 1681620392
transform 1 0 1308 0 1 2375
box -3 -3 3 3
use BUFX2  BUFX2_1
timestamp 1681620392
transform -1 0 1304 0 1 2370
box -5 -3 28 105
use FILL  FILL_244
timestamp 1681620392
transform 1 0 1304 0 1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_21
timestamp 1681620392
transform 1 0 1312 0 1 2370
box -8 -3 32 105
use M3_M2  M3_M2_944
timestamp 1681620392
transform 1 0 1404 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_70
timestamp 1681620392
transform 1 0 1336 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_71
timestamp 1681620392
transform 1 0 1432 0 1 2370
box -8 -3 104 105
use NAND2X1  NAND2X1_48
timestamp 1681620392
transform 1 0 1528 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_49
timestamp 1681620392
transform 1 0 1552 0 1 2370
box -8 -3 32 105
use OAI21X1  OAI21X1_80
timestamp 1681620392
transform 1 0 1576 0 1 2370
box -8 -3 34 105
use NAND2X1  NAND2X1_50
timestamp 1681620392
transform 1 0 1608 0 1 2370
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_72
timestamp 1681620392
transform 1 0 1632 0 1 2370
box -8 -3 104 105
use NAND2X1  NAND2X1_51
timestamp 1681620392
transform -1 0 1752 0 1 2370
box -8 -3 32 105
use BUFX2  BUFX2_2
timestamp 1681620392
transform -1 0 1776 0 1 2370
box -5 -3 28 105
use BUFX2  BUFX2_3
timestamp 1681620392
transform -1 0 1800 0 1 2370
box -5 -3 28 105
use NAND2X1  NAND2X1_52
timestamp 1681620392
transform 1 0 1800 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_53
timestamp 1681620392
transform -1 0 1848 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_54
timestamp 1681620392
transform -1 0 1872 0 1 2370
box -8 -3 32 105
use OAI21X1  OAI21X1_81
timestamp 1681620392
transform -1 0 1904 0 1 2370
box -8 -3 34 105
use M3_M2  M3_M2_945
timestamp 1681620392
transform 1 0 1996 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_73
timestamp 1681620392
transform 1 0 1904 0 1 2370
box -8 -3 104 105
use NAND2X1  NAND2X1_55
timestamp 1681620392
transform 1 0 2000 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_56
timestamp 1681620392
transform 1 0 2024 0 1 2370
box -8 -3 32 105
use OAI21X1  OAI21X1_82
timestamp 1681620392
transform 1 0 2048 0 1 2370
box -8 -3 34 105
use M3_M2  M3_M2_946
timestamp 1681620392
transform 1 0 2092 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_74
timestamp 1681620392
transform -1 0 2176 0 1 2370
box -8 -3 104 105
use M3_M2  M3_M2_947
timestamp 1681620392
transform 1 0 2196 0 1 2375
box -3 -3 3 3
use OAI21X1  OAI21X1_83
timestamp 1681620392
transform 1 0 2176 0 1 2370
box -8 -3 34 105
use NAND2X1  NAND2X1_57
timestamp 1681620392
transform 1 0 2208 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_58
timestamp 1681620392
transform 1 0 2232 0 1 2370
box -8 -3 32 105
use M3_M2  M3_M2_948
timestamp 1681620392
transform 1 0 2292 0 1 2375
box -3 -3 3 3
use BUFX2  BUFX2_4
timestamp 1681620392
transform 1 0 2256 0 1 2370
box -5 -3 28 105
use FILL  FILL_245
timestamp 1681620392
transform 1 0 2280 0 1 2370
box -8 -3 16 105
use FILL  FILL_246
timestamp 1681620392
transform 1 0 2288 0 1 2370
box -8 -3 16 105
use NAND2X1  NAND2X1_59
timestamp 1681620392
transform 1 0 2296 0 1 2370
box -8 -3 32 105
use FILL  FILL_247
timestamp 1681620392
transform 1 0 2320 0 1 2370
box -8 -3 16 105
use FILL  FILL_248
timestamp 1681620392
transform 1 0 2328 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_84
timestamp 1681620392
transform -1 0 2368 0 1 2370
box -8 -3 34 105
use FILL  FILL_249
timestamp 1681620392
transform 1 0 2368 0 1 2370
box -8 -3 16 105
use FILL  FILL_250
timestamp 1681620392
transform 1 0 2376 0 1 2370
box -8 -3 16 105
use NAND2X1  NAND2X1_63
timestamp 1681620392
transform 1 0 2384 0 1 2370
box -8 -3 32 105
use FILL  FILL_265
timestamp 1681620392
transform 1 0 2408 0 1 2370
box -8 -3 16 105
use FILL  FILL_266
timestamp 1681620392
transform 1 0 2416 0 1 2370
box -8 -3 16 105
use FILL  FILL_269
timestamp 1681620392
transform 1 0 2424 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_86
timestamp 1681620392
transform -1 0 2464 0 1 2370
box -8 -3 34 105
use NAND2X1  NAND2X1_65
timestamp 1681620392
transform -1 0 2488 0 1 2370
box -8 -3 32 105
use FILL  FILL_270
timestamp 1681620392
transform 1 0 2488 0 1 2370
box -8 -3 16 105
use FILL  FILL_274
timestamp 1681620392
transform 1 0 2496 0 1 2370
box -8 -3 16 105
use FILL  FILL_276
timestamp 1681620392
transform 1 0 2504 0 1 2370
box -8 -3 16 105
use FILL  FILL_278
timestamp 1681620392
transform 1 0 2512 0 1 2370
box -8 -3 16 105
use FILL  FILL_279
timestamp 1681620392
transform 1 0 2520 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_87
timestamp 1681620392
transform -1 0 2560 0 1 2370
box -8 -3 34 105
use M3_M2  M3_M2_949
timestamp 1681620392
transform 1 0 2572 0 1 2375
box -3 -3 3 3
use FILL  FILL_280
timestamp 1681620392
transform 1 0 2560 0 1 2370
box -8 -3 16 105
use NAND2X1  NAND2X1_68
timestamp 1681620392
transform -1 0 2592 0 1 2370
box -8 -3 32 105
use FILL  FILL_281
timestamp 1681620392
transform 1 0 2592 0 1 2370
box -8 -3 16 105
use FILL  FILL_282
timestamp 1681620392
transform 1 0 2600 0 1 2370
box -8 -3 16 105
use FILL  FILL_283
timestamp 1681620392
transform 1 0 2608 0 1 2370
box -8 -3 16 105
use FILL  FILL_284
timestamp 1681620392
transform 1 0 2616 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_82
timestamp 1681620392
transform 1 0 2624 0 1 2370
box -9 -3 26 105
use FILL  FILL_285
timestamp 1681620392
transform 1 0 2640 0 1 2370
box -8 -3 16 105
use AND2X2  AND2X2_7
timestamp 1681620392
transform -1 0 2680 0 1 2370
box -8 -3 40 105
use FILL  FILL_286
timestamp 1681620392
transform 1 0 2680 0 1 2370
box -8 -3 16 105
use FILL  FILL_287
timestamp 1681620392
transform 1 0 2688 0 1 2370
box -8 -3 16 105
use FILL  FILL_288
timestamp 1681620392
transform 1 0 2696 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_950
timestamp 1681620392
transform 1 0 2716 0 1 2375
box -3 -3 3 3
use FILL  FILL_289
timestamp 1681620392
transform 1 0 2704 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_88
timestamp 1681620392
transform -1 0 2744 0 1 2370
box -8 -3 34 105
use INVX2  INVX2_83
timestamp 1681620392
transform 1 0 2744 0 1 2370
box -9 -3 26 105
use FILL  FILL_290
timestamp 1681620392
transform 1 0 2760 0 1 2370
box -8 -3 16 105
use FILL  FILL_291
timestamp 1681620392
transform 1 0 2768 0 1 2370
box -8 -3 16 105
use FILL  FILL_292
timestamp 1681620392
transform 1 0 2776 0 1 2370
box -8 -3 16 105
use FILL  FILL_293
timestamp 1681620392
transform 1 0 2784 0 1 2370
box -8 -3 16 105
use FILL  FILL_294
timestamp 1681620392
transform 1 0 2792 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_89
timestamp 1681620392
transform 1 0 2800 0 1 2370
box -8 -3 34 105
use NAND2X1  NAND2X1_69
timestamp 1681620392
transform -1 0 2856 0 1 2370
box -8 -3 32 105
use FILL  FILL_295
timestamp 1681620392
transform 1 0 2856 0 1 2370
box -8 -3 16 105
use FILL  FILL_296
timestamp 1681620392
transform 1 0 2864 0 1 2370
box -8 -3 16 105
use FILL  FILL_297
timestamp 1681620392
transform 1 0 2872 0 1 2370
box -8 -3 16 105
use FILL  FILL_298
timestamp 1681620392
transform 1 0 2880 0 1 2370
box -8 -3 16 105
use FILL  FILL_299
timestamp 1681620392
transform 1 0 2888 0 1 2370
box -8 -3 16 105
use NAND2X1  NAND2X1_70
timestamp 1681620392
transform -1 0 2920 0 1 2370
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_85
timestamp 1681620392
transform 1 0 2920 0 1 2370
box -8 -3 104 105
use Project_Top_VIA0  Project_Top_VIA0_13
timestamp 1681620392
transform 1 0 3043 0 1 2370
box -10 -3 10 3
use M3_M2  M3_M2_951
timestamp 1681620392
transform 1 0 68 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_966
timestamp 1681620392
transform 1 0 68 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_1159
timestamp 1681620392
transform 1 0 68 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_1164
timestamp 1681620392
transform 1 0 68 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_1063
timestamp 1681620392
transform 1 0 68 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_1165
timestamp 1681620392
transform 1 0 92 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1166
timestamp 1681620392
transform 1 0 116 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1221
timestamp 1681620392
transform 1 0 116 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1167
timestamp 1681620392
transform 1 0 132 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1222
timestamp 1681620392
transform 1 0 132 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1223
timestamp 1681620392
transform 1 0 148 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1301
timestamp 1681620392
transform 1 0 132 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_1039
timestamp 1681620392
transform 1 0 132 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_967
timestamp 1681620392
transform 1 0 172 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_1168
timestamp 1681620392
transform 1 0 164 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1169
timestamp 1681620392
transform 1 0 172 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1224
timestamp 1681620392
transform 1 0 180 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1302
timestamp 1681620392
transform 1 0 188 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_1004
timestamp 1681620392
transform 1 0 204 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_1225
timestamp 1681620392
transform 1 0 212 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_952
timestamp 1681620392
transform 1 0 260 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_953
timestamp 1681620392
transform 1 0 276 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_973
timestamp 1681620392
transform 1 0 244 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_1170
timestamp 1681620392
transform 1 0 276 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1171
timestamp 1681620392
transform 1 0 292 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_1005
timestamp 1681620392
transform 1 0 236 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1006
timestamp 1681620392
transform 1 0 260 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_1303
timestamp 1681620392
transform 1 0 212 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_1040
timestamp 1681620392
transform 1 0 196 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1021
timestamp 1681620392
transform 1 0 220 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_1304
timestamp 1681620392
transform 1 0 236 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1305
timestamp 1681620392
transform 1 0 252 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1306
timestamp 1681620392
transform 1 0 260 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1330
timestamp 1681620392
transform 1 0 204 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_1331
timestamp 1681620392
transform 1 0 244 0 1 2305
box -2 -2 2 2
use M3_M2  M3_M2_1007
timestamp 1681620392
transform 1 0 284 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_1226
timestamp 1681620392
transform 1 0 292 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1307
timestamp 1681620392
transform 1 0 284 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1332
timestamp 1681620392
transform 1 0 268 0 1 2305
box -2 -2 2 2
use M3_M2  M3_M2_974
timestamp 1681620392
transform 1 0 324 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_1172
timestamp 1681620392
transform 1 0 324 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1173
timestamp 1681620392
transform 1 0 332 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1227
timestamp 1681620392
transform 1 0 316 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1228
timestamp 1681620392
transform 1 0 324 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1229
timestamp 1681620392
transform 1 0 340 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_1022
timestamp 1681620392
transform 1 0 324 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_975
timestamp 1681620392
transform 1 0 364 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_1308
timestamp 1681620392
transform 1 0 356 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_1041
timestamp 1681620392
transform 1 0 356 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_976
timestamp 1681620392
transform 1 0 396 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_1174
timestamp 1681620392
transform 1 0 388 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1175
timestamp 1681620392
transform 1 0 404 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1230
timestamp 1681620392
transform 1 0 388 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1231
timestamp 1681620392
transform 1 0 404 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1232
timestamp 1681620392
transform 1 0 412 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1309
timestamp 1681620392
transform 1 0 372 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1310
timestamp 1681620392
transform 1 0 396 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_1023
timestamp 1681620392
transform 1 0 404 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_1333
timestamp 1681620392
transform 1 0 380 0 1 2305
box -2 -2 2 2
use M3_M2  M3_M2_1042
timestamp 1681620392
transform 1 0 388 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1064
timestamp 1681620392
transform 1 0 404 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_1311
timestamp 1681620392
transform 1 0 420 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_1043
timestamp 1681620392
transform 1 0 420 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_1176
timestamp 1681620392
transform 1 0 444 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_1008
timestamp 1681620392
transform 1 0 444 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_1233
timestamp 1681620392
transform 1 0 452 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1234
timestamp 1681620392
transform 1 0 460 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_1024
timestamp 1681620392
transform 1 0 452 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_1312
timestamp 1681620392
transform 1 0 468 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_1065
timestamp 1681620392
transform 1 0 460 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1025
timestamp 1681620392
transform 1 0 476 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_977
timestamp 1681620392
transform 1 0 500 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_1235
timestamp 1681620392
transform 1 0 500 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1313
timestamp 1681620392
transform 1 0 492 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1314
timestamp 1681620392
transform 1 0 516 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1315
timestamp 1681620392
transform 1 0 540 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1177
timestamp 1681620392
transform 1 0 548 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_1066
timestamp 1681620392
transform 1 0 540 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_998
timestamp 1681620392
transform 1 0 556 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_1178
timestamp 1681620392
transform 1 0 572 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1179
timestamp 1681620392
transform 1 0 588 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_999
timestamp 1681620392
transform 1 0 612 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_978
timestamp 1681620392
transform 1 0 700 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_1160
timestamp 1681620392
transform 1 0 708 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_1180
timestamp 1681620392
transform 1 0 692 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1181
timestamp 1681620392
transform 1 0 700 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1236
timestamp 1681620392
transform 1 0 572 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1237
timestamp 1681620392
transform 1 0 612 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1238
timestamp 1681620392
transform 1 0 668 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1239
timestamp 1681620392
transform 1 0 676 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1240
timestamp 1681620392
transform 1 0 684 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_1026
timestamp 1681620392
transform 1 0 572 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1027
timestamp 1681620392
transform 1 0 676 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1028
timestamp 1681620392
transform 1 0 692 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1044
timestamp 1681620392
transform 1 0 668 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_979
timestamp 1681620392
transform 1 0 724 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_1182
timestamp 1681620392
transform 1 0 724 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1241
timestamp 1681620392
transform 1 0 748 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_980
timestamp 1681620392
transform 1 0 812 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1000
timestamp 1681620392
transform 1 0 820 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_1242
timestamp 1681620392
transform 1 0 812 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1243
timestamp 1681620392
transform 1 0 820 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1183
timestamp 1681620392
transform 1 0 836 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_1009
timestamp 1681620392
transform 1 0 828 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_1184
timestamp 1681620392
transform 1 0 852 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1161
timestamp 1681620392
transform 1 0 868 0 1 2345
box -2 -2 2 2
use M3_M2  M3_M2_1001
timestamp 1681620392
transform 1 0 868 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_1244
timestamp 1681620392
transform 1 0 860 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1245
timestamp 1681620392
transform 1 0 868 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1185
timestamp 1681620392
transform 1 0 892 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1246
timestamp 1681620392
transform 1 0 884 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1247
timestamp 1681620392
transform 1 0 908 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_1010
timestamp 1681620392
transform 1 0 916 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_1316
timestamp 1681620392
transform 1 0 900 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1334
timestamp 1681620392
transform 1 0 892 0 1 2305
box -2 -2 2 2
use M3_M2  M3_M2_981
timestamp 1681620392
transform 1 0 940 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_1186
timestamp 1681620392
transform 1 0 940 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1317
timestamp 1681620392
transform 1 0 932 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_954
timestamp 1681620392
transform 1 0 1036 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_982
timestamp 1681620392
transform 1 0 1020 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_1187
timestamp 1681620392
transform 1 0 1020 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1681620392
transform 1 0 1028 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1248
timestamp 1681620392
transform 1 0 948 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1249
timestamp 1681620392
transform 1 0 964 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1250
timestamp 1681620392
transform 1 0 988 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1318
timestamp 1681620392
transform 1 0 972 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_1045
timestamp 1681620392
transform 1 0 948 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1011
timestamp 1681620392
transform 1 0 996 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_983
timestamp 1681620392
transform 1 0 1068 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_1189
timestamp 1681620392
transform 1 0 1060 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1251
timestamp 1681620392
transform 1 0 1028 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1252
timestamp 1681620392
transform 1 0 1044 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1681620392
transform 1 0 996 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1320
timestamp 1681620392
transform 1 0 1004 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1321
timestamp 1681620392
transform 1 0 1020 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1335
timestamp 1681620392
transform 1 0 980 0 1 2305
box -2 -2 2 2
use M3_M2  M3_M2_1046
timestamp 1681620392
transform 1 0 1004 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1067
timestamp 1681620392
transform 1 0 988 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1012
timestamp 1681620392
transform 1 0 1060 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_968
timestamp 1681620392
transform 1 0 1084 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_1253
timestamp 1681620392
transform 1 0 1076 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1322
timestamp 1681620392
transform 1 0 1076 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_1068
timestamp 1681620392
transform 1 0 1076 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_969
timestamp 1681620392
transform 1 0 1100 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_970
timestamp 1681620392
transform 1 0 1204 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_1190
timestamp 1681620392
transform 1 0 1116 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1191
timestamp 1681620392
transform 1 0 1204 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_971
timestamp 1681620392
transform 1 0 1236 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_1162
timestamp 1681620392
transform 1 0 1236 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_1192
timestamp 1681620392
transform 1 0 1228 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1193
timestamp 1681620392
transform 1 0 1244 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1254
timestamp 1681620392
transform 1 0 1108 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1255
timestamp 1681620392
transform 1 0 1124 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1256
timestamp 1681620392
transform 1 0 1180 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1257
timestamp 1681620392
transform 1 0 1220 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_1029
timestamp 1681620392
transform 1 0 1116 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1047
timestamp 1681620392
transform 1 0 1124 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1075
timestamp 1681620392
transform 1 0 1108 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1013
timestamp 1681620392
transform 1 0 1228 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_1258
timestamp 1681620392
transform 1 0 1236 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_1014
timestamp 1681620392
transform 1 0 1244 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1030
timestamp 1681620392
transform 1 0 1220 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_1259
timestamp 1681620392
transform 1 0 1260 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_1069
timestamp 1681620392
transform 1 0 1252 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_955
timestamp 1681620392
transform 1 0 1300 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_984
timestamp 1681620392
transform 1 0 1292 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_1163
timestamp 1681620392
transform 1 0 1300 0 1 2345
box -2 -2 2 2
use M3_M2  M3_M2_972
timestamp 1681620392
transform 1 0 1316 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_1194
timestamp 1681620392
transform 1 0 1300 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1681620392
transform 1 0 1308 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_1031
timestamp 1681620392
transform 1 0 1300 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_985
timestamp 1681620392
transform 1 0 1388 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_956
timestamp 1681620392
transform 1 0 1428 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_1196
timestamp 1681620392
transform 1 0 1404 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1197
timestamp 1681620392
transform 1 0 1420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1260
timestamp 1681620392
transform 1 0 1316 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1261
timestamp 1681620392
transform 1 0 1324 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1262
timestamp 1681620392
transform 1 0 1372 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_1032
timestamp 1681620392
transform 1 0 1324 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1070
timestamp 1681620392
transform 1 0 1316 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1076
timestamp 1681620392
transform 1 0 1308 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1048
timestamp 1681620392
transform 1 0 1428 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_1263
timestamp 1681620392
transform 1 0 1444 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_1049
timestamp 1681620392
transform 1 0 1444 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_1198
timestamp 1681620392
transform 1 0 1468 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_1002
timestamp 1681620392
transform 1 0 1540 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1003
timestamp 1681620392
transform 1 0 1556 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_1264
timestamp 1681620392
transform 1 0 1492 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1265
timestamp 1681620392
transform 1 0 1548 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1266
timestamp 1681620392
transform 1 0 1556 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1199
timestamp 1681620392
transform 1 0 1564 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_1015
timestamp 1681620392
transform 1 0 1564 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_957
timestamp 1681620392
transform 1 0 1588 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_958
timestamp 1681620392
transform 1 0 1612 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_1200
timestamp 1681620392
transform 1 0 1668 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1267
timestamp 1681620392
transform 1 0 1580 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1268
timestamp 1681620392
transform 1 0 1588 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1269
timestamp 1681620392
transform 1 0 1620 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_1033
timestamp 1681620392
transform 1 0 1596 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1034
timestamp 1681620392
transform 1 0 1620 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1016
timestamp 1681620392
transform 1 0 1684 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_1323
timestamp 1681620392
transform 1 0 1684 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_986
timestamp 1681620392
transform 1 0 1748 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_987
timestamp 1681620392
transform 1 0 1804 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_988
timestamp 1681620392
transform 1 0 1828 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_1201
timestamp 1681620392
transform 1 0 1716 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1202
timestamp 1681620392
transform 1 0 1732 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1203
timestamp 1681620392
transform 1 0 1820 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1270
timestamp 1681620392
transform 1 0 1708 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1271
timestamp 1681620392
transform 1 0 1764 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1272
timestamp 1681620392
transform 1 0 1812 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_1035
timestamp 1681620392
transform 1 0 1732 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1036
timestamp 1681620392
transform 1 0 1780 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1050
timestamp 1681620392
transform 1 0 1820 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_959
timestamp 1681620392
transform 1 0 1972 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_989
timestamp 1681620392
transform 1 0 1868 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_990
timestamp 1681620392
transform 1 0 1884 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_1204
timestamp 1681620392
transform 1 0 1860 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_960
timestamp 1681620392
transform 1 0 2004 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_991
timestamp 1681620392
transform 1 0 1980 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_992
timestamp 1681620392
transform 1 0 2060 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_1205
timestamp 1681620392
transform 1 0 1884 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1206
timestamp 1681620392
transform 1 0 1900 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1273
timestamp 1681620392
transform 1 0 1844 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1274
timestamp 1681620392
transform 1 0 1868 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1207
timestamp 1681620392
transform 1 0 1996 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_961
timestamp 1681620392
transform 1 0 2132 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_1208
timestamp 1681620392
transform 1 0 2092 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1275
timestamp 1681620392
transform 1 0 1932 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1276
timestamp 1681620392
transform 1 0 1980 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1277
timestamp 1681620392
transform 1 0 2044 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1278
timestamp 1681620392
transform 1 0 2076 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1279
timestamp 1681620392
transform 1 0 2140 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1280
timestamp 1681620392
transform 1 0 2172 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_1051
timestamp 1681620392
transform 1 0 1900 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1052
timestamp 1681620392
transform 1 0 1996 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1053
timestamp 1681620392
transform 1 0 2044 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1054
timestamp 1681620392
transform 1 0 2092 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1077
timestamp 1681620392
transform 1 0 2052 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1078
timestamp 1681620392
transform 1 0 2076 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1079
timestamp 1681620392
transform 1 0 2100 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_962
timestamp 1681620392
transform 1 0 2284 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_993
timestamp 1681620392
transform 1 0 2212 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_1209
timestamp 1681620392
transform 1 0 2196 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1210
timestamp 1681620392
transform 1 0 2292 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1281
timestamp 1681620392
transform 1 0 2236 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1282
timestamp 1681620392
transform 1 0 2276 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1283
timestamp 1681620392
transform 1 0 2316 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1284
timestamp 1681620392
transform 1 0 2372 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_1055
timestamp 1681620392
transform 1 0 2340 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1056
timestamp 1681620392
transform 1 0 2372 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_1324
timestamp 1681620392
transform 1 0 2412 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_1071
timestamp 1681620392
transform 1 0 2412 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_1285
timestamp 1681620392
transform 1 0 2428 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1286
timestamp 1681620392
transform 1 0 2436 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1211
timestamp 1681620392
transform 1 0 2468 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1287
timestamp 1681620392
transform 1 0 2460 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1325
timestamp 1681620392
transform 1 0 2460 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1212
timestamp 1681620392
transform 1 0 2484 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1681620392
transform 1 0 2484 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_1057
timestamp 1681620392
transform 1 0 2460 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1058
timestamp 1681620392
transform 1 0 2476 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1072
timestamp 1681620392
transform 1 0 2484 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_1288
timestamp 1681620392
transform 1 0 2500 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1213
timestamp 1681620392
transform 1 0 2556 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1289
timestamp 1681620392
transform 1 0 2548 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1214
timestamp 1681620392
transform 1 0 2580 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1290
timestamp 1681620392
transform 1 0 2572 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1327
timestamp 1681620392
transform 1 0 2572 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_1073
timestamp 1681620392
transform 1 0 2572 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_963
timestamp 1681620392
transform 1 0 2692 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_964
timestamp 1681620392
transform 1 0 2748 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_994
timestamp 1681620392
transform 1 0 2660 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_1215
timestamp 1681620392
transform 1 0 2612 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_995
timestamp 1681620392
transform 1 0 2708 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_996
timestamp 1681620392
transform 1 0 2740 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_1216
timestamp 1681620392
transform 1 0 2708 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1291
timestamp 1681620392
transform 1 0 2596 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1292
timestamp 1681620392
transform 1 0 2660 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1293
timestamp 1681620392
transform 1 0 2692 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1328
timestamp 1681620392
transform 1 0 2596 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_1037
timestamp 1681620392
transform 1 0 2636 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1038
timestamp 1681620392
transform 1 0 2660 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1074
timestamp 1681620392
transform 1 0 2596 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1017
timestamp 1681620392
transform 1 0 2708 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_965
timestamp 1681620392
transform 1 0 2884 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_997
timestamp 1681620392
transform 1 0 2900 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_1217
timestamp 1681620392
transform 1 0 2804 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1218
timestamp 1681620392
transform 1 0 2892 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1294
timestamp 1681620392
transform 1 0 2732 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1295
timestamp 1681620392
transform 1 0 2788 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_1059
timestamp 1681620392
transform 1 0 2700 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1060
timestamp 1681620392
transform 1 0 2732 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1018
timestamp 1681620392
transform 1 0 2804 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_1296
timestamp 1681620392
transform 1 0 2828 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_1019
timestamp 1681620392
transform 1 0 2836 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_1219
timestamp 1681620392
transform 1 0 2916 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1220
timestamp 1681620392
transform 1 0 2932 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1297
timestamp 1681620392
transform 1 0 2884 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1298
timestamp 1681620392
transform 1 0 2900 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_1061
timestamp 1681620392
transform 1 0 2876 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1020
timestamp 1681620392
transform 1 0 2932 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_1299
timestamp 1681620392
transform 1 0 2956 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1300
timestamp 1681620392
transform 1 0 3012 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1329
timestamp 1681620392
transform 1 0 2916 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_1062
timestamp 1681620392
transform 1 0 2916 0 1 2305
box -3 -3 3 3
use Project_Top_VIA0  Project_Top_VIA0_14
timestamp 1681620392
transform 1 0 24 0 1 2270
box -10 -3 10 3
use FILL  FILL_214
timestamp 1681620392
transform 1 0 72 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_1080
timestamp 1681620392
transform 1 0 116 0 1 2275
box -3 -3 3 3
use OR2X1  OR2X1_2
timestamp 1681620392
transform 1 0 80 0 -1 2370
box -8 -3 40 105
use INVX2  INVX2_67
timestamp 1681620392
transform 1 0 112 0 -1 2370
box -9 -3 26 105
use OAI21X1  OAI21X1_75
timestamp 1681620392
transform -1 0 160 0 -1 2370
box -8 -3 34 105
use FILL  FILL_215
timestamp 1681620392
transform 1 0 160 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_68
timestamp 1681620392
transform 1 0 168 0 -1 2370
box -9 -3 26 105
use FILL  FILL_216
timestamp 1681620392
transform 1 0 184 0 -1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_22
timestamp 1681620392
transform -1 0 224 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_23
timestamp 1681620392
transform 1 0 224 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_24
timestamp 1681620392
transform -1 0 288 0 -1 2370
box -8 -3 40 105
use INVX2  INVX2_69
timestamp 1681620392
transform 1 0 288 0 -1 2370
box -9 -3 26 105
use FILL  FILL_217
timestamp 1681620392
transform 1 0 304 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_70
timestamp 1681620392
transform -1 0 328 0 -1 2370
box -9 -3 26 105
use NAND2X1  NAND2X1_43
timestamp 1681620392
transform 1 0 328 0 -1 2370
box -8 -3 32 105
use FILL  FILL_218
timestamp 1681620392
transform 1 0 352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_219
timestamp 1681620392
transform 1 0 360 0 -1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_25
timestamp 1681620392
transform -1 0 400 0 -1 2370
box -8 -3 40 105
use NAND2X1  NAND2X1_44
timestamp 1681620392
transform 1 0 400 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_45
timestamp 1681620392
transform -1 0 448 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_46
timestamp 1681620392
transform 1 0 448 0 -1 2370
box -8 -3 32 105
use FILL  FILL_220
timestamp 1681620392
transform 1 0 472 0 -1 2370
box -8 -3 16 105
use FILL  FILL_229
timestamp 1681620392
transform 1 0 480 0 -1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_27
timestamp 1681620392
transform 1 0 488 0 -1 2370
box -8 -3 40 105
use FILL  FILL_230
timestamp 1681620392
transform 1 0 520 0 -1 2370
box -8 -3 16 105
use FILL  FILL_231
timestamp 1681620392
transform 1 0 528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_232
timestamp 1681620392
transform 1 0 536 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_77
timestamp 1681620392
transform -1 0 576 0 -1 2370
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_67
timestamp 1681620392
transform 1 0 576 0 -1 2370
box -8 -3 104 105
use M3_M2  M3_M2_1081
timestamp 1681620392
transform 1 0 684 0 1 2275
box -3 -3 3 3
use INVX2  INVX2_72
timestamp 1681620392
transform -1 0 688 0 -1 2370
box -9 -3 26 105
use NOR2X1  NOR2X1_19
timestamp 1681620392
transform -1 0 712 0 -1 2370
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_68
timestamp 1681620392
transform 1 0 712 0 -1 2370
box -8 -3 104 105
use FILL  FILL_233
timestamp 1681620392
transform 1 0 808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_251
timestamp 1681620392
transform 1 0 816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_252
timestamp 1681620392
transform 1 0 824 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_76
timestamp 1681620392
transform 1 0 832 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_77
timestamp 1681620392
transform 1 0 848 0 -1 2370
box -9 -3 26 105
use NOR2X1  NOR2X1_22
timestamp 1681620392
transform 1 0 864 0 -1 2370
box -8 -3 32 105
use FILL  FILL_253
timestamp 1681620392
transform 1 0 888 0 -1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_30
timestamp 1681620392
transform 1 0 896 0 -1 2370
box -8 -3 40 105
use FILL  FILL_254
timestamp 1681620392
transform 1 0 928 0 -1 2370
box -8 -3 16 105
use AND2X2  AND2X2_5
timestamp 1681620392
transform 1 0 936 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_31
timestamp 1681620392
transform -1 0 1000 0 -1 2370
box -8 -3 40 105
use NAND2X1  NAND2X1_60
timestamp 1681620392
transform -1 0 1024 0 -1 2370
box -8 -3 32 105
use OAI21X1  OAI21X1_85
timestamp 1681620392
transform -1 0 1056 0 -1 2370
box -8 -3 34 105
use NAND2X1  NAND2X1_61
timestamp 1681620392
transform 1 0 1056 0 -1 2370
box -8 -3 32 105
use FILL  FILL_255
timestamp 1681620392
transform 1 0 1080 0 -1 2370
box -8 -3 16 105
use AND2X2  AND2X2_6
timestamp 1681620392
transform -1 0 1120 0 -1 2370
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_75
timestamp 1681620392
transform -1 0 1216 0 -1 2370
box -8 -3 104 105
use NOR2X1  NOR2X1_23
timestamp 1681620392
transform -1 0 1240 0 -1 2370
box -8 -3 32 105
use INVX2  INVX2_78
timestamp 1681620392
transform 1 0 1240 0 -1 2370
box -9 -3 26 105
use FILL  FILL_256
timestamp 1681620392
transform 1 0 1256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_257
timestamp 1681620392
transform 1 0 1264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_258
timestamp 1681620392
transform 1 0 1272 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_79
timestamp 1681620392
transform -1 0 1296 0 -1 2370
box -9 -3 26 105
use NOR2X1  NOR2X1_24
timestamp 1681620392
transform 1 0 1296 0 -1 2370
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_76
timestamp 1681620392
transform -1 0 1416 0 -1 2370
box -8 -3 104 105
use BUFX2  BUFX2_5
timestamp 1681620392
transform -1 0 1440 0 -1 2370
box -5 -3 28 105
use FILL  FILL_259
timestamp 1681620392
transform 1 0 1440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_260
timestamp 1681620392
transform 1 0 1448 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_77
timestamp 1681620392
transform 1 0 1456 0 -1 2370
box -8 -3 104 105
use INVX2  INVX2_80
timestamp 1681620392
transform -1 0 1568 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_81
timestamp 1681620392
transform 1 0 1568 0 -1 2370
box -9 -3 26 105
use M3_M2  M3_M2_1082
timestamp 1681620392
transform 1 0 1636 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1083
timestamp 1681620392
transform 1 0 1668 0 1 2275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_78
timestamp 1681620392
transform -1 0 1680 0 -1 2370
box -8 -3 104 105
use FILL  FILL_261
timestamp 1681620392
transform 1 0 1680 0 -1 2370
box -8 -3 16 105
use FILL  FILL_262
timestamp 1681620392
transform 1 0 1688 0 -1 2370
box -8 -3 16 105
use NAND2X1  NAND2X1_62
timestamp 1681620392
transform -1 0 1720 0 -1 2370
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_79
timestamp 1681620392
transform 1 0 1720 0 -1 2370
box -8 -3 104 105
use BUFX2  BUFX2_6
timestamp 1681620392
transform -1 0 1840 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_7
timestamp 1681620392
transform 1 0 1840 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_8
timestamp 1681620392
transform 1 0 1864 0 -1 2370
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_80
timestamp 1681620392
transform 1 0 1888 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_81
timestamp 1681620392
transform 1 0 1984 0 -1 2370
box -8 -3 104 105
use M3_M2  M3_M2_1084
timestamp 1681620392
transform 1 0 2140 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1085
timestamp 1681620392
transform 1 0 2172 0 1 2275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_82
timestamp 1681620392
transform 1 0 2080 0 -1 2370
box -8 -3 104 105
use FILL  FILL_263
timestamp 1681620392
transform 1 0 2176 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_83
timestamp 1681620392
transform 1 0 2184 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_84
timestamp 1681620392
transform 1 0 2280 0 -1 2370
box -8 -3 104 105
use FILL  FILL_264
timestamp 1681620392
transform 1 0 2376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_267
timestamp 1681620392
transform 1 0 2384 0 -1 2370
box -8 -3 16 105
use NAND2X1  NAND2X1_64
timestamp 1681620392
transform 1 0 2392 0 -1 2370
box -8 -3 32 105
use FILL  FILL_268
timestamp 1681620392
transform 1 0 2416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_271
timestamp 1681620392
transform 1 0 2424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_272
timestamp 1681620392
transform 1 0 2432 0 -1 2370
box -8 -3 16 105
use NAND2X1  NAND2X1_66
timestamp 1681620392
transform 1 0 2440 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_67
timestamp 1681620392
transform 1 0 2464 0 -1 2370
box -8 -3 32 105
use FILL  FILL_273
timestamp 1681620392
transform 1 0 2488 0 -1 2370
box -8 -3 16 105
use FILL  FILL_275
timestamp 1681620392
transform 1 0 2496 0 -1 2370
box -8 -3 16 105
use FILL  FILL_277
timestamp 1681620392
transform 1 0 2504 0 -1 2370
box -8 -3 16 105
use FILL  FILL_300
timestamp 1681620392
transform 1 0 2512 0 -1 2370
box -8 -3 16 105
use BUFX2  BUFX2_9
timestamp 1681620392
transform -1 0 2544 0 -1 2370
box -5 -3 28 105
use FILL  FILL_301
timestamp 1681620392
transform 1 0 2544 0 -1 2370
box -8 -3 16 105
use NAND2X1  NAND2X1_71
timestamp 1681620392
transform 1 0 2552 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_72
timestamp 1681620392
transform 1 0 2576 0 -1 2370
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_86
timestamp 1681620392
transform 1 0 2600 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_87
timestamp 1681620392
transform 1 0 2696 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_88
timestamp 1681620392
transform 1 0 2792 0 -1 2370
box -8 -3 104 105
use OAI21X1  OAI21X1_90
timestamp 1681620392
transform 1 0 2888 0 -1 2370
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_89
timestamp 1681620392
transform 1 0 2920 0 -1 2370
box -8 -3 104 105
use Project_Top_VIA0  Project_Top_VIA0_15
timestamp 1681620392
transform 1 0 3067 0 1 2270
box -10 -3 10 3
use M2_M1  M2_M1_1382
timestamp 1681620392
transform 1 0 68 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1383
timestamp 1681620392
transform 1 0 124 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1466
timestamp 1681620392
transform 1 0 156 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1199
timestamp 1681620392
transform 1 0 156 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1091
timestamp 1681620392
transform 1 0 276 0 1 2255
box -3 -3 3 3
use M2_M1  M2_M1_1384
timestamp 1681620392
transform 1 0 236 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1385
timestamp 1681620392
transform 1 0 276 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1467
timestamp 1681620392
transform 1 0 188 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1200
timestamp 1681620392
transform 1 0 188 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1201
timestamp 1681620392
transform 1 0 236 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1099
timestamp 1681620392
transform 1 0 292 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_1343
timestamp 1681620392
transform 1 0 292 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1386
timestamp 1681620392
transform 1 0 292 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1387
timestamp 1681620392
transform 1 0 308 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1388
timestamp 1681620392
transform 1 0 316 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1468
timestamp 1681620392
transform 1 0 292 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1202
timestamp 1681620392
transform 1 0 292 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1086
timestamp 1681620392
transform 1 0 332 0 1 2265
box -3 -3 3 3
use M2_M1  M2_M1_1336
timestamp 1681620392
transform 1 0 348 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_1344
timestamp 1681620392
transform 1 0 332 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1469
timestamp 1681620392
transform 1 0 324 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1203
timestamp 1681620392
transform 1 0 324 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1134
timestamp 1681620392
transform 1 0 348 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1087
timestamp 1681620392
transform 1 0 372 0 1 2265
box -3 -3 3 3
use M2_M1  M2_M1_1345
timestamp 1681620392
transform 1 0 356 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1389
timestamp 1681620392
transform 1 0 340 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1390
timestamp 1681620392
transform 1 0 364 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1544
timestamp 1681620392
transform 1 0 364 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_1237
timestamp 1681620392
transform 1 0 340 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1113
timestamp 1681620392
transform 1 0 380 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1135
timestamp 1681620392
transform 1 0 388 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1100
timestamp 1681620392
transform 1 0 420 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1101
timestamp 1681620392
transform 1 0 468 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1102
timestamp 1681620392
transform 1 0 484 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_1337
timestamp 1681620392
transform 1 0 436 0 1 2235
box -2 -2 2 2
use M3_M2  M3_M2_1114
timestamp 1681620392
transform 1 0 444 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_1346
timestamp 1681620392
transform 1 0 420 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1391
timestamp 1681620392
transform 1 0 380 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1392
timestamp 1681620392
transform 1 0 388 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1393
timestamp 1681620392
transform 1 0 404 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1136
timestamp 1681620392
transform 1 0 428 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_1347
timestamp 1681620392
transform 1 0 444 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1348
timestamp 1681620392
transform 1 0 476 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1394
timestamp 1681620392
transform 1 0 428 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1395
timestamp 1681620392
transform 1 0 452 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1396
timestamp 1681620392
transform 1 0 468 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1470
timestamp 1681620392
transform 1 0 412 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1471
timestamp 1681620392
transform 1 0 476 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1472
timestamp 1681620392
transform 1 0 484 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1204
timestamp 1681620392
transform 1 0 452 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1205
timestamp 1681620392
transform 1 0 484 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1137
timestamp 1681620392
transform 1 0 516 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_1349
timestamp 1681620392
transform 1 0 628 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1397
timestamp 1681620392
transform 1 0 532 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1398
timestamp 1681620392
transform 1 0 564 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1473
timestamp 1681620392
transform 1 0 508 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1474
timestamp 1681620392
transform 1 0 524 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1190
timestamp 1681620392
transform 1 0 532 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1157
timestamp 1681620392
transform 1 0 628 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1475
timestamp 1681620392
transform 1 0 612 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1476
timestamp 1681620392
transform 1 0 628 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1206
timestamp 1681620392
transform 1 0 564 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1207
timestamp 1681620392
transform 1 0 612 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1088
timestamp 1681620392
transform 1 0 700 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1103
timestamp 1681620392
transform 1 0 708 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1104
timestamp 1681620392
transform 1 0 756 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1105
timestamp 1681620392
transform 1 0 780 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1106
timestamp 1681620392
transform 1 0 796 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1138
timestamp 1681620392
transform 1 0 684 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_1350
timestamp 1681620392
transform 1 0 700 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_1139
timestamp 1681620392
transform 1 0 804 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_1399
timestamp 1681620392
transform 1 0 684 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1477
timestamp 1681620392
transform 1 0 652 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1478
timestamp 1681620392
transform 1 0 668 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1479
timestamp 1681620392
transform 1 0 676 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1158
timestamp 1681620392
transform 1 0 700 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1400
timestamp 1681620392
transform 1 0 740 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1159
timestamp 1681620392
transform 1 0 748 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1401
timestamp 1681620392
transform 1 0 796 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1402
timestamp 1681620392
transform 1 0 804 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1403
timestamp 1681620392
transform 1 0 812 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1480
timestamp 1681620392
transform 1 0 700 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1481
timestamp 1681620392
transform 1 0 716 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1191
timestamp 1681620392
transform 1 0 796 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1208
timestamp 1681620392
transform 1 0 716 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1238
timestamp 1681620392
transform 1 0 788 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_1351
timestamp 1681620392
transform 1 0 828 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_1115
timestamp 1681620392
transform 1 0 844 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_1338
timestamp 1681620392
transform 1 0 868 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_1352
timestamp 1681620392
transform 1 0 852 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1404
timestamp 1681620392
transform 1 0 836 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1209
timestamp 1681620392
transform 1 0 828 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1140
timestamp 1681620392
transform 1 0 868 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_1482
timestamp 1681620392
transform 1 0 844 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1239
timestamp 1681620392
transform 1 0 868 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_1353
timestamp 1681620392
transform 1 0 884 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_1160
timestamp 1681620392
transform 1 0 884 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1483
timestamp 1681620392
transform 1 0 884 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1141
timestamp 1681620392
transform 1 0 908 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_1405
timestamp 1681620392
transform 1 0 900 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1406
timestamp 1681620392
transform 1 0 908 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1192
timestamp 1681620392
transform 1 0 900 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_1484
timestamp 1681620392
transform 1 0 908 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1116
timestamp 1681620392
transform 1 0 924 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_1354
timestamp 1681620392
transform 1 0 924 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_1161
timestamp 1681620392
transform 1 0 924 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1162
timestamp 1681620392
transform 1 0 940 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1407
timestamp 1681620392
transform 1 0 948 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1485
timestamp 1681620392
transform 1 0 924 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1486
timestamp 1681620392
transform 1 0 948 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1210
timestamp 1681620392
transform 1 0 948 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1117
timestamp 1681620392
transform 1 0 988 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_1355
timestamp 1681620392
transform 1 0 980 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1408
timestamp 1681620392
transform 1 0 972 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1163
timestamp 1681620392
transform 1 0 980 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1142
timestamp 1681620392
transform 1 0 1012 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_1409
timestamp 1681620392
transform 1 0 988 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1193
timestamp 1681620392
transform 1 0 972 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_1487
timestamp 1681620392
transform 1 0 980 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1164
timestamp 1681620392
transform 1 0 1004 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1118
timestamp 1681620392
transform 1 0 1028 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_1410
timestamp 1681620392
transform 1 0 1012 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1411
timestamp 1681620392
transform 1 0 1020 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1488
timestamp 1681620392
transform 1 0 1012 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1545
timestamp 1681620392
transform 1 0 1028 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_1092
timestamp 1681620392
transform 1 0 1076 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1119
timestamp 1681620392
transform 1 0 1060 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_1339
timestamp 1681620392
transform 1 0 1068 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_1340
timestamp 1681620392
transform 1 0 1092 0 1 2235
box -2 -2 2 2
use M3_M2  M3_M2_1143
timestamp 1681620392
transform 1 0 1052 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_1356
timestamp 1681620392
transform 1 0 1060 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_1144
timestamp 1681620392
transform 1 0 1092 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_1412
timestamp 1681620392
transform 1 0 1052 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1413
timestamp 1681620392
transform 1 0 1076 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1414
timestamp 1681620392
transform 1 0 1092 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1489
timestamp 1681620392
transform 1 0 1052 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1357
timestamp 1681620392
transform 1 0 1108 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_1145
timestamp 1681620392
transform 1 0 1124 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_1415
timestamp 1681620392
transform 1 0 1116 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1416
timestamp 1681620392
transform 1 0 1124 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1490
timestamp 1681620392
transform 1 0 1108 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1240
timestamp 1681620392
transform 1 0 1116 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1093
timestamp 1681620392
transform 1 0 1164 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1120
timestamp 1681620392
transform 1 0 1164 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_1417
timestamp 1681620392
transform 1 0 1164 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1418
timestamp 1681620392
transform 1 0 1180 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1491
timestamp 1681620392
transform 1 0 1140 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1211
timestamp 1681620392
transform 1 0 1140 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_1358
timestamp 1681620392
transform 1 0 1228 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_1165
timestamp 1681620392
transform 1 0 1204 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1419
timestamp 1681620392
transform 1 0 1228 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1492
timestamp 1681620392
transform 1 0 1172 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1493
timestamp 1681620392
transform 1 0 1196 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1494
timestamp 1681620392
transform 1 0 1212 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1212
timestamp 1681620392
transform 1 0 1196 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1194
timestamp 1681620392
transform 1 0 1220 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_1546
timestamp 1681620392
transform 1 0 1204 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_1241
timestamp 1681620392
transform 1 0 1172 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1213
timestamp 1681620392
transform 1 0 1228 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_1359
timestamp 1681620392
transform 1 0 1244 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1420
timestamp 1681620392
transform 1 0 1252 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1495
timestamp 1681620392
transform 1 0 1244 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1146
timestamp 1681620392
transform 1 0 1268 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1094
timestamp 1681620392
transform 1 0 1348 0 1 2255
box -3 -3 3 3
use M2_M1  M2_M1_1341
timestamp 1681620392
transform 1 0 1292 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_1342
timestamp 1681620392
transform 1 0 1300 0 1 2235
box -2 -2 2 2
use M3_M2  M3_M2_1121
timestamp 1681620392
transform 1 0 1308 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1122
timestamp 1681620392
transform 1 0 1324 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_1360
timestamp 1681620392
transform 1 0 1276 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_1147
timestamp 1681620392
transform 1 0 1300 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_1361
timestamp 1681620392
transform 1 0 1308 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1362
timestamp 1681620392
transform 1 0 1316 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1421
timestamp 1681620392
transform 1 0 1268 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1166
timestamp 1681620392
transform 1 0 1276 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1422
timestamp 1681620392
transform 1 0 1300 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1496
timestamp 1681620392
transform 1 0 1276 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1214
timestamp 1681620392
transform 1 0 1276 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1148
timestamp 1681620392
transform 1 0 1324 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_1363
timestamp 1681620392
transform 1 0 1340 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1364
timestamp 1681620392
transform 1 0 1348 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_1149
timestamp 1681620392
transform 1 0 1364 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_1365
timestamp 1681620392
transform 1 0 1380 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1423
timestamp 1681620392
transform 1 0 1324 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1167
timestamp 1681620392
transform 1 0 1340 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1150
timestamp 1681620392
transform 1 0 1396 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_1424
timestamp 1681620392
transform 1 0 1364 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1425
timestamp 1681620392
transform 1 0 1372 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1168
timestamp 1681620392
transform 1 0 1380 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1426
timestamp 1681620392
transform 1 0 1396 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1497
timestamp 1681620392
transform 1 0 1348 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1498
timestamp 1681620392
transform 1 0 1372 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1499
timestamp 1681620392
transform 1 0 1404 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1500
timestamp 1681620392
transform 1 0 1412 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1215
timestamp 1681620392
transform 1 0 1372 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1216
timestamp 1681620392
transform 1 0 1404 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1242
timestamp 1681620392
transform 1 0 1396 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_1427
timestamp 1681620392
transform 1 0 1428 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1501
timestamp 1681620392
transform 1 0 1436 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1217
timestamp 1681620392
transform 1 0 1436 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1095
timestamp 1681620392
transform 1 0 1460 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1107
timestamp 1681620392
transform 1 0 1452 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_1366
timestamp 1681620392
transform 1 0 1452 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1428
timestamp 1681620392
transform 1 0 1460 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1108
timestamp 1681620392
transform 1 0 1500 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1123
timestamp 1681620392
transform 1 0 1484 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1151
timestamp 1681620392
transform 1 0 1476 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1124
timestamp 1681620392
transform 1 0 1508 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_1367
timestamp 1681620392
transform 1 0 1500 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1368
timestamp 1681620392
transform 1 0 1508 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1429
timestamp 1681620392
transform 1 0 1484 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1169
timestamp 1681620392
transform 1 0 1492 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1430
timestamp 1681620392
transform 1 0 1500 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1170
timestamp 1681620392
transform 1 0 1508 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1431
timestamp 1681620392
transform 1 0 1524 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1502
timestamp 1681620392
transform 1 0 1476 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1503
timestamp 1681620392
transform 1 0 1484 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1218
timestamp 1681620392
transform 1 0 1484 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_1504
timestamp 1681620392
transform 1 0 1508 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1505
timestamp 1681620392
transform 1 0 1532 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1219
timestamp 1681620392
transform 1 0 1516 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1220
timestamp 1681620392
transform 1 0 1532 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1152
timestamp 1681620392
transform 1 0 1548 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1109
timestamp 1681620392
transform 1 0 1564 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_1369
timestamp 1681620392
transform 1 0 1564 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1432
timestamp 1681620392
transform 1 0 1612 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1506
timestamp 1681620392
transform 1 0 1588 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1507
timestamp 1681620392
transform 1 0 1596 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1110
timestamp 1681620392
transform 1 0 1740 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_1370
timestamp 1681620392
transform 1 0 1740 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1433
timestamp 1681620392
transform 1 0 1660 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1434
timestamp 1681620392
transform 1 0 1716 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1435
timestamp 1681620392
transform 1 0 1732 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1508
timestamp 1681620392
transform 1 0 1620 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1509
timestamp 1681620392
transform 1 0 1636 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1221
timestamp 1681620392
transform 1 0 1620 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1243
timestamp 1681620392
transform 1 0 1724 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1171
timestamp 1681620392
transform 1 0 1748 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1436
timestamp 1681620392
transform 1 0 1756 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1172
timestamp 1681620392
transform 1 0 1764 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1173
timestamp 1681620392
transform 1 0 1780 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1437
timestamp 1681620392
transform 1 0 1820 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1438
timestamp 1681620392
transform 1 0 1860 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1174
timestamp 1681620392
transform 1 0 1868 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1439
timestamp 1681620392
transform 1 0 1884 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1510
timestamp 1681620392
transform 1 0 1764 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1511
timestamp 1681620392
transform 1 0 1780 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1512
timestamp 1681620392
transform 1 0 1868 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1222
timestamp 1681620392
transform 1 0 1764 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1223
timestamp 1681620392
transform 1 0 1812 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1244
timestamp 1681620392
transform 1 0 1772 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1125
timestamp 1681620392
transform 1 0 1940 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_1371
timestamp 1681620392
transform 1 0 1940 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1440
timestamp 1681620392
transform 1 0 1924 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1111
timestamp 1681620392
transform 1 0 2052 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1126
timestamp 1681620392
transform 1 0 2052 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_1372
timestamp 1681620392
transform 1 0 2044 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1441
timestamp 1681620392
transform 1 0 1988 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1175
timestamp 1681620392
transform 1 0 2004 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1442
timestamp 1681620392
transform 1 0 2036 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1176
timestamp 1681620392
transform 1 0 2044 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1443
timestamp 1681620392
transform 1 0 2052 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1513
timestamp 1681620392
transform 1 0 1908 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1514
timestamp 1681620392
transform 1 0 1916 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1515
timestamp 1681620392
transform 1 0 1940 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1516
timestamp 1681620392
transform 1 0 1956 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1224
timestamp 1681620392
transform 1 0 1916 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1225
timestamp 1681620392
transform 1 0 1932 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_1444
timestamp 1681620392
transform 1 0 2076 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1517
timestamp 1681620392
transform 1 0 2060 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1518
timestamp 1681620392
transform 1 0 2068 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1226
timestamp 1681620392
transform 1 0 2068 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1096
timestamp 1681620392
transform 1 0 2124 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1127
timestamp 1681620392
transform 1 0 2124 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_1373
timestamp 1681620392
transform 1 0 2116 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1374
timestamp 1681620392
transform 1 0 2124 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_1177
timestamp 1681620392
transform 1 0 2108 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1445
timestamp 1681620392
transform 1 0 2116 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1519
timestamp 1681620392
transform 1 0 2092 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1520
timestamp 1681620392
transform 1 0 2100 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1128
timestamp 1681620392
transform 1 0 2180 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_1375
timestamp 1681620392
transform 1 0 2180 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1446
timestamp 1681620392
transform 1 0 2164 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1521
timestamp 1681620392
transform 1 0 2140 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1522
timestamp 1681620392
transform 1 0 2148 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1523
timestamp 1681620392
transform 1 0 2172 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1245
timestamp 1681620392
transform 1 0 2172 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_1447
timestamp 1681620392
transform 1 0 2204 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1524
timestamp 1681620392
transform 1 0 2196 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1227
timestamp 1681620392
transform 1 0 2196 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_1376
timestamp 1681620392
transform 1 0 2244 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1448
timestamp 1681620392
transform 1 0 2220 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1525
timestamp 1681620392
transform 1 0 2212 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1246
timestamp 1681620392
transform 1 0 2212 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1178
timestamp 1681620392
transform 1 0 2244 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1526
timestamp 1681620392
transform 1 0 2236 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1195
timestamp 1681620392
transform 1 0 2260 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_1449
timestamp 1681620392
transform 1 0 2276 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1450
timestamp 1681620392
transform 1 0 2284 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1527
timestamp 1681620392
transform 1 0 2268 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1528
timestamp 1681620392
transform 1 0 2292 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1377
timestamp 1681620392
transform 1 0 2324 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_1179
timestamp 1681620392
transform 1 0 2324 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1529
timestamp 1681620392
transform 1 0 2316 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1228
timestamp 1681620392
transform 1 0 2316 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1097
timestamp 1681620392
transform 1 0 2428 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1180
timestamp 1681620392
transform 1 0 2356 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1098
timestamp 1681620392
transform 1 0 2460 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1129
timestamp 1681620392
transform 1 0 2516 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1130
timestamp 1681620392
transform 1 0 2540 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_1378
timestamp 1681620392
transform 1 0 2540 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1451
timestamp 1681620392
transform 1 0 2380 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1452
timestamp 1681620392
transform 1 0 2436 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1530
timestamp 1681620392
transform 1 0 2340 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1531
timestamp 1681620392
transform 1 0 2356 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1229
timestamp 1681620392
transform 1 0 2388 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1181
timestamp 1681620392
transform 1 0 2452 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1453
timestamp 1681620392
transform 1 0 2484 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1454
timestamp 1681620392
transform 1 0 2532 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1455
timestamp 1681620392
transform 1 0 2540 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1532
timestamp 1681620392
transform 1 0 2452 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1230
timestamp 1681620392
transform 1 0 2452 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1182
timestamp 1681620392
transform 1 0 2564 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1533
timestamp 1681620392
transform 1 0 2564 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1231
timestamp 1681620392
transform 1 0 2564 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1153
timestamp 1681620392
transform 1 0 2580 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1131
timestamp 1681620392
transform 1 0 2612 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_1379
timestamp 1681620392
transform 1 0 2596 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1456
timestamp 1681620392
transform 1 0 2580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1457
timestamp 1681620392
transform 1 0 2588 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1183
timestamp 1681620392
transform 1 0 2604 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1184
timestamp 1681620392
transform 1 0 2620 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1154
timestamp 1681620392
transform 1 0 2636 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_1534
timestamp 1681620392
transform 1 0 2628 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1458
timestamp 1681620392
transform 1 0 2644 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1459
timestamp 1681620392
transform 1 0 2652 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1535
timestamp 1681620392
transform 1 0 2644 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1196
timestamp 1681620392
transform 1 0 2652 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1089
timestamp 1681620392
transform 1 0 2668 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1155
timestamp 1681620392
transform 1 0 2668 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1112
timestamp 1681620392
transform 1 0 2708 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_1380
timestamp 1681620392
transform 1 0 2708 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_1132
timestamp 1681620392
transform 1 0 2740 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1156
timestamp 1681620392
transform 1 0 2804 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1185
timestamp 1681620392
transform 1 0 2676 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1460
timestamp 1681620392
transform 1 0 2684 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1186
timestamp 1681620392
transform 1 0 2692 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1187
timestamp 1681620392
transform 1 0 2708 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1188
timestamp 1681620392
transform 1 0 2724 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1461
timestamp 1681620392
transform 1 0 2780 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_1189
timestamp 1681620392
transform 1 0 2788 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_1462
timestamp 1681620392
transform 1 0 2820 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1463
timestamp 1681620392
transform 1 0 2860 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1464
timestamp 1681620392
transform 1 0 2916 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1465
timestamp 1681620392
transform 1 0 2932 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1536
timestamp 1681620392
transform 1 0 2668 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1232
timestamp 1681620392
transform 1 0 2660 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1197
timestamp 1681620392
transform 1 0 2692 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_1537
timestamp 1681620392
transform 1 0 2700 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1547
timestamp 1681620392
transform 1 0 2668 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_1198
timestamp 1681620392
transform 1 0 2716 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_1538
timestamp 1681620392
transform 1 0 2724 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1539
timestamp 1681620392
transform 1 0 2740 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1233
timestamp 1681620392
transform 1 0 2724 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_1540
timestamp 1681620392
transform 1 0 2836 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1541
timestamp 1681620392
transform 1 0 2924 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1234
timestamp 1681620392
transform 1 0 2836 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1235
timestamp 1681620392
transform 1 0 2868 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1236
timestamp 1681620392
transform 1 0 2924 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1247
timestamp 1681620392
transform 1 0 2924 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_1542
timestamp 1681620392
transform 1 0 2956 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_1133
timestamp 1681620392
transform 1 0 2972 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_1381
timestamp 1681620392
transform 1 0 2972 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_1090
timestamp 1681620392
transform 1 0 3012 0 1 2265
box -3 -3 3 3
use M2_M1  M2_M1_1543
timestamp 1681620392
transform 1 0 3012 0 1 2205
box -2 -2 2 2
use Project_Top_VIA0  Project_Top_VIA0_16
timestamp 1681620392
transform 1 0 48 0 1 2170
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_90
timestamp 1681620392
transform -1 0 168 0 1 2170
box -8 -3 104 105
use FILL  FILL_302
timestamp 1681620392
transform 1 0 168 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_91
timestamp 1681620392
transform 1 0 176 0 1 2170
box -8 -3 104 105
use INVX2  INVX2_84
timestamp 1681620392
transform 1 0 272 0 1 2170
box -9 -3 26 105
use OAI21X1  OAI21X1_91
timestamp 1681620392
transform -1 0 320 0 1 2170
box -8 -3 34 105
use FILL  FILL_303
timestamp 1681620392
transform 1 0 320 0 1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_32
timestamp 1681620392
transform 1 0 328 0 1 2170
box -8 -3 40 105
use NOR2X1  NOR2X1_25
timestamp 1681620392
transform 1 0 360 0 1 2170
box -8 -3 32 105
use AND2X2  AND2X2_8
timestamp 1681620392
transform -1 0 416 0 1 2170
box -8 -3 40 105
use M3_M2  M3_M2_1248
timestamp 1681620392
transform 1 0 452 0 1 2175
box -3 -3 3 3
use NAND3X1  NAND3X1_33
timestamp 1681620392
transform 1 0 416 0 1 2170
box -8 -3 40 105
use AND2X2  AND2X2_9
timestamp 1681620392
transform -1 0 480 0 1 2170
box -8 -3 40 105
use M3_M2  M3_M2_1249
timestamp 1681620392
transform 1 0 508 0 1 2175
box -3 -3 3 3
use OAI21X1  OAI21X1_92
timestamp 1681620392
transform -1 0 512 0 1 2170
box -8 -3 34 105
use INVX2  INVX2_85
timestamp 1681620392
transform -1 0 528 0 1 2170
box -9 -3 26 105
use M3_M2  M3_M2_1250
timestamp 1681620392
transform 1 0 572 0 1 2175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_92
timestamp 1681620392
transform -1 0 624 0 1 2170
box -8 -3 104 105
use M3_M2  M3_M2_1251
timestamp 1681620392
transform 1 0 652 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1252
timestamp 1681620392
transform 1 0 676 0 1 2175
box -3 -3 3 3
use OAI21X1  OAI21X1_93
timestamp 1681620392
transform -1 0 656 0 1 2170
box -8 -3 34 105
use INVX2  INVX2_86
timestamp 1681620392
transform -1 0 672 0 1 2170
box -9 -3 26 105
use M3_M2  M3_M2_1253
timestamp 1681620392
transform 1 0 716 0 1 2175
box -3 -3 3 3
use OAI21X1  OAI21X1_94
timestamp 1681620392
transform 1 0 672 0 1 2170
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_98
timestamp 1681620392
transform 1 0 704 0 1 2170
box -8 -3 104 105
use INVX2  INVX2_88
timestamp 1681620392
transform -1 0 816 0 1 2170
box -9 -3 26 105
use FILL  FILL_305
timestamp 1681620392
transform 1 0 816 0 1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_74
timestamp 1681620392
transform -1 0 848 0 1 2170
box -8 -3 32 105
use NAND3X1  NAND3X1_34
timestamp 1681620392
transform 1 0 848 0 1 2170
box -8 -3 40 105
use FILL  FILL_306
timestamp 1681620392
transform 1 0 880 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_89
timestamp 1681620392
transform 1 0 888 0 1 2170
box -9 -3 26 105
use NAND2X1  NAND2X1_75
timestamp 1681620392
transform 1 0 904 0 1 2170
box -8 -3 32 105
use INVX2  INVX2_93
timestamp 1681620392
transform 1 0 928 0 1 2170
box -9 -3 26 105
use FILL  FILL_313
timestamp 1681620392
transform 1 0 944 0 1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_79
timestamp 1681620392
transform 1 0 952 0 1 2170
box -8 -3 32 105
use AND2X2  AND2X2_10
timestamp 1681620392
transform 1 0 976 0 1 2170
box -8 -3 40 105
use INVX2  INVX2_94
timestamp 1681620392
transform 1 0 1008 0 1 2170
box -9 -3 26 105
use FILL  FILL_317
timestamp 1681620392
transform 1 0 1024 0 1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_27
timestamp 1681620392
transform 1 0 1032 0 1 2170
box -8 -3 32 105
use NAND3X1  NAND3X1_35
timestamp 1681620392
transform -1 0 1088 0 1 2170
box -8 -3 40 105
use NAND2X1  NAND2X1_80
timestamp 1681620392
transform 1 0 1088 0 1 2170
box -8 -3 32 105
use OAI21X1  OAI21X1_98
timestamp 1681620392
transform 1 0 1112 0 1 2170
box -8 -3 34 105
use AND2X2  AND2X2_11
timestamp 1681620392
transform -1 0 1176 0 1 2170
box -8 -3 40 105
use OR2X1  OR2X1_4
timestamp 1681620392
transform -1 0 1208 0 1 2170
box -8 -3 40 105
use INVX2  INVX2_95
timestamp 1681620392
transform 1 0 1208 0 1 2170
box -9 -3 26 105
use NAND2X1  NAND2X1_81
timestamp 1681620392
transform -1 0 1248 0 1 2170
box -8 -3 32 105
use FILL  FILL_318
timestamp 1681620392
transform 1 0 1248 0 1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_82
timestamp 1681620392
transform -1 0 1280 0 1 2170
box -8 -3 32 105
use NAND3X1  NAND3X1_36
timestamp 1681620392
transform -1 0 1312 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_37
timestamp 1681620392
transform 1 0 1312 0 1 2170
box -8 -3 40 105
use OAI21X1  OAI21X1_99
timestamp 1681620392
transform -1 0 1376 0 1 2170
box -8 -3 34 105
use M3_M2  M3_M2_1254
timestamp 1681620392
transform 1 0 1412 0 1 2175
box -3 -3 3 3
use OAI21X1  OAI21X1_100
timestamp 1681620392
transform -1 0 1408 0 1 2170
box -8 -3 34 105
use BUFX2  BUFX2_10
timestamp 1681620392
transform -1 0 1432 0 1 2170
box -5 -3 28 105
use INVX2  INVX2_96
timestamp 1681620392
transform 1 0 1432 0 1 2170
box -9 -3 26 105
use FILL  FILL_319
timestamp 1681620392
transform 1 0 1448 0 1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_83
timestamp 1681620392
transform -1 0 1480 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_84
timestamp 1681620392
transform 1 0 1480 0 1 2170
box -8 -3 32 105
use OAI21X1  OAI21X1_101
timestamp 1681620392
transform -1 0 1536 0 1 2170
box -8 -3 34 105
use FILL  FILL_320
timestamp 1681620392
transform 1 0 1536 0 1 2170
box -8 -3 16 105
use FILL  FILL_321
timestamp 1681620392
transform 1 0 1544 0 1 2170
box -8 -3 16 105
use FILL  FILL_322
timestamp 1681620392
transform 1 0 1552 0 1 2170
box -8 -3 16 105
use FILL  FILL_323
timestamp 1681620392
transform 1 0 1560 0 1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_85
timestamp 1681620392
transform -1 0 1592 0 1 2170
box -8 -3 32 105
use OAI21X1  OAI21X1_102
timestamp 1681620392
transform -1 0 1624 0 1 2170
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_99
timestamp 1681620392
transform 1 0 1624 0 1 2170
box -8 -3 104 105
use NAND2X1  NAND2X1_86
timestamp 1681620392
transform 1 0 1720 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_87
timestamp 1681620392
transform -1 0 1768 0 1 2170
box -8 -3 32 105
use M3_M2  M3_M2_1255
timestamp 1681620392
transform 1 0 1828 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1256
timestamp 1681620392
transform 1 0 1860 0 1 2175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_100
timestamp 1681620392
transform 1 0 1768 0 1 2170
box -8 -3 104 105
use BUFX2  BUFX2_11
timestamp 1681620392
transform -1 0 1888 0 1 2170
box -5 -3 28 105
use BUFX2  BUFX2_12
timestamp 1681620392
transform 1 0 1888 0 1 2170
box -5 -3 28 105
use OAI21X1  OAI21X1_103
timestamp 1681620392
transform 1 0 1912 0 1 2170
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_101
timestamp 1681620392
transform 1 0 1944 0 1 2170
box -8 -3 104 105
use NAND2X1  NAND2X1_88
timestamp 1681620392
transform -1 0 2064 0 1 2170
box -8 -3 32 105
use OAI21X1  OAI21X1_104
timestamp 1681620392
transform 1 0 2064 0 1 2170
box -8 -3 34 105
use NAND2X1  NAND2X1_89
timestamp 1681620392
transform 1 0 2096 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_90
timestamp 1681620392
transform -1 0 2144 0 1 2170
box -8 -3 32 105
use OAI21X1  OAI21X1_105
timestamp 1681620392
transform -1 0 2176 0 1 2170
box -8 -3 34 105
use NAND2X1  NAND2X1_91
timestamp 1681620392
transform -1 0 2200 0 1 2170
box -8 -3 32 105
use FILL  FILL_324
timestamp 1681620392
transform 1 0 2200 0 1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_114
timestamp 1681620392
transform 1 0 2208 0 1 2170
box -8 -3 34 105
use NAND2X1  NAND2X1_98
timestamp 1681620392
transform -1 0 2264 0 1 2170
box -8 -3 32 105
use FILL  FILL_341
timestamp 1681620392
transform 1 0 2264 0 1 2170
box -8 -3 16 105
use FILL  FILL_342
timestamp 1681620392
transform 1 0 2272 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_1257
timestamp 1681620392
transform 1 0 2292 0 1 2175
box -3 -3 3 3
use FILL  FILL_343
timestamp 1681620392
transform 1 0 2280 0 1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_115
timestamp 1681620392
transform 1 0 2288 0 1 2170
box -8 -3 34 105
use M3_M2  M3_M2_1258
timestamp 1681620392
transform 1 0 2332 0 1 2175
box -3 -3 3 3
use NAND2X1  NAND2X1_99
timestamp 1681620392
transform -1 0 2344 0 1 2170
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_107
timestamp 1681620392
transform 1 0 2344 0 1 2170
box -8 -3 104 105
use M3_M2  M3_M2_1259
timestamp 1681620392
transform 1 0 2460 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1260
timestamp 1681620392
transform 1 0 2492 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1261
timestamp 1681620392
transform 1 0 2532 0 1 2175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_108
timestamp 1681620392
transform 1 0 2440 0 1 2170
box -8 -3 104 105
use NAND2X1  NAND2X1_100
timestamp 1681620392
transform -1 0 2560 0 1 2170
box -8 -3 32 105
use FILL  FILL_344
timestamp 1681620392
transform 1 0 2560 0 1 2170
box -8 -3 16 105
use FILL  FILL_345
timestamp 1681620392
transform 1 0 2568 0 1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_101
timestamp 1681620392
transform 1 0 2576 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_102
timestamp 1681620392
transform -1 0 2624 0 1 2170
box -8 -3 32 105
use FILL  FILL_346
timestamp 1681620392
transform 1 0 2624 0 1 2170
box -8 -3 16 105
use FILL  FILL_347
timestamp 1681620392
transform 1 0 2632 0 1 2170
box -8 -3 16 105
use FILL  FILL_348
timestamp 1681620392
transform 1 0 2640 0 1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_29
timestamp 1681620392
transform -1 0 2672 0 1 2170
box -8 -3 32 105
use OAI21X1  OAI21X1_116
timestamp 1681620392
transform 1 0 2672 0 1 2170
box -8 -3 34 105
use NAND2X1  NAND2X1_103
timestamp 1681620392
transform -1 0 2728 0 1 2170
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_109
timestamp 1681620392
transform 1 0 2728 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_110
timestamp 1681620392
transform 1 0 2824 0 1 2170
box -8 -3 104 105
use OAI21X1  OAI21X1_117
timestamp 1681620392
transform 1 0 2920 0 1 2170
box -8 -3 34 105
use FILL  FILL_349
timestamp 1681620392
transform 1 0 2952 0 1 2170
box -8 -3 16 105
use FILL  FILL_350
timestamp 1681620392
transform 1 0 2960 0 1 2170
box -8 -3 16 105
use FILL  FILL_351
timestamp 1681620392
transform 1 0 2968 0 1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_104
timestamp 1681620392
transform -1 0 3000 0 1 2170
box -8 -3 32 105
use FILL  FILL_352
timestamp 1681620392
transform 1 0 3000 0 1 2170
box -8 -3 16 105
use FILL  FILL_353
timestamp 1681620392
transform 1 0 3008 0 1 2170
box -8 -3 16 105
use Project_Top_VIA0  Project_Top_VIA0_17
timestamp 1681620392
transform 1 0 3043 0 1 2170
box -10 -3 10 3
use M2_M1  M2_M1_1551
timestamp 1681620392
transform 1 0 84 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1552
timestamp 1681620392
transform 1 0 172 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1635
timestamp 1681620392
transform 1 0 124 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1636
timestamp 1681620392
transform 1 0 164 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1371
timestamp 1681620392
transform 1 0 172 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1343
timestamp 1681620392
transform 1 0 188 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_1553
timestamp 1681620392
transform 1 0 204 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1554
timestamp 1681620392
transform 1 0 228 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_1344
timestamp 1681620392
transform 1 0 268 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_1555
timestamp 1681620392
transform 1 0 316 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1637
timestamp 1681620392
transform 1 0 188 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1638
timestamp 1681620392
transform 1 0 196 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1639
timestamp 1681620392
transform 1 0 212 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1640
timestamp 1681620392
transform 1 0 228 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1641
timestamp 1681620392
transform 1 0 236 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1642
timestamp 1681620392
transform 1 0 268 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1709
timestamp 1681620392
transform 1 0 188 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1372
timestamp 1681620392
transform 1 0 212 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1310
timestamp 1681620392
transform 1 0 388 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1311
timestamp 1681620392
transform 1 0 428 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1556
timestamp 1681620392
transform 1 0 340 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_1345
timestamp 1681620392
transform 1 0 420 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_1557
timestamp 1681620392
transform 1 0 428 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1643
timestamp 1681620392
transform 1 0 388 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1644
timestamp 1681620392
transform 1 0 420 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1710
timestamp 1681620392
transform 1 0 428 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1262
timestamp 1681620392
transform 1 0 468 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_1558
timestamp 1681620392
transform 1 0 452 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_1346
timestamp 1681620392
transform 1 0 460 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_1559
timestamp 1681620392
transform 1 0 468 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1560
timestamp 1681620392
transform 1 0 564 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1645
timestamp 1681620392
transform 1 0 484 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1646
timestamp 1681620392
transform 1 0 524 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1283
timestamp 1681620392
transform 1 0 668 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1312
timestamp 1681620392
transform 1 0 588 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1313
timestamp 1681620392
transform 1 0 612 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1561
timestamp 1681620392
transform 1 0 588 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1562
timestamp 1681620392
transform 1 0 676 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1647
timestamp 1681620392
transform 1 0 628 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1356
timestamp 1681620392
transform 1 0 660 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1263
timestamp 1681620392
transform 1 0 708 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_1648
timestamp 1681620392
transform 1 0 668 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1649
timestamp 1681620392
transform 1 0 684 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1650
timestamp 1681620392
transform 1 0 700 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1711
timestamp 1681620392
transform 1 0 708 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1563
timestamp 1681620392
transform 1 0 724 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_1357
timestamp 1681620392
transform 1 0 732 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1264
timestamp 1681620392
transform 1 0 748 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1314
timestamp 1681620392
transform 1 0 740 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1564
timestamp 1681620392
transform 1 0 740 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1565
timestamp 1681620392
transform 1 0 748 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1651
timestamp 1681620392
transform 1 0 740 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1373
timestamp 1681620392
transform 1 0 740 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1347
timestamp 1681620392
transform 1 0 756 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_1566
timestamp 1681620392
transform 1 0 764 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1652
timestamp 1681620392
transform 1 0 764 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1374
timestamp 1681620392
transform 1 0 764 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1414
timestamp 1681620392
transform 1 0 772 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1265
timestamp 1681620392
transform 1 0 804 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1315
timestamp 1681620392
transform 1 0 796 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1548
timestamp 1681620392
transform 1 0 804 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1567
timestamp 1681620392
transform 1 0 820 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1712
timestamp 1681620392
transform 1 0 812 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1316
timestamp 1681620392
transform 1 0 844 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1568
timestamp 1681620392
transform 1 0 844 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_1358
timestamp 1681620392
transform 1 0 828 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_1653
timestamp 1681620392
transform 1 0 836 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1359
timestamp 1681620392
transform 1 0 844 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1284
timestamp 1681620392
transform 1 0 860 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_1569
timestamp 1681620392
transform 1 0 860 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1570
timestamp 1681620392
transform 1 0 876 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1571
timestamp 1681620392
transform 1 0 884 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1654
timestamp 1681620392
transform 1 0 852 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1655
timestamp 1681620392
transform 1 0 868 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1385
timestamp 1681620392
transform 1 0 820 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1406
timestamp 1681620392
transform 1 0 812 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_1713
timestamp 1681620392
transform 1 0 844 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1407
timestamp 1681620392
transform 1 0 868 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1266
timestamp 1681620392
transform 1 0 908 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_1572
timestamp 1681620392
transform 1 0 900 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1656
timestamp 1681620392
transform 1 0 908 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1375
timestamp 1681620392
transform 1 0 892 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_1714
timestamp 1681620392
transform 1 0 900 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1376
timestamp 1681620392
transform 1 0 908 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1386
timestamp 1681620392
transform 1 0 900 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_1657
timestamp 1681620392
transform 1 0 924 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1285
timestamp 1681620392
transform 1 0 956 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_1573
timestamp 1681620392
transform 1 0 956 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_1267
timestamp 1681620392
transform 1 0 980 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_1574
timestamp 1681620392
transform 1 0 980 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1658
timestamp 1681620392
transform 1 0 980 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1360
timestamp 1681620392
transform 1 0 988 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1268
timestamp 1681620392
transform 1 0 1108 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1286
timestamp 1681620392
transform 1 0 1020 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1287
timestamp 1681620392
transform 1 0 1084 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1317
timestamp 1681620392
transform 1 0 1044 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1575
timestamp 1681620392
transform 1 0 1020 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1659
timestamp 1681620392
transform 1 0 996 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1715
timestamp 1681620392
transform 1 0 964 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1377
timestamp 1681620392
transform 1 0 972 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_1716
timestamp 1681620392
transform 1 0 988 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1361
timestamp 1681620392
transform 1 0 1004 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1269
timestamp 1681620392
transform 1 0 1140 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_1576
timestamp 1681620392
transform 1 0 1148 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1577
timestamp 1681620392
transform 1 0 1156 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1660
timestamp 1681620392
transform 1 0 1044 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1661
timestamp 1681620392
transform 1 0 1100 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1662
timestamp 1681620392
transform 1 0 1116 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1717
timestamp 1681620392
transform 1 0 1004 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1387
timestamp 1681620392
transform 1 0 996 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1408
timestamp 1681620392
transform 1 0 980 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1362
timestamp 1681620392
transform 1 0 1124 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_1663
timestamp 1681620392
transform 1 0 1140 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1718
timestamp 1681620392
transform 1 0 1108 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1378
timestamp 1681620392
transform 1 0 1116 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_1719
timestamp 1681620392
transform 1 0 1132 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1388
timestamp 1681620392
transform 1 0 1108 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_1739
timestamp 1681620392
transform 1 0 1124 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_1409
timestamp 1681620392
transform 1 0 1116 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1389
timestamp 1681620392
transform 1 0 1156 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1318
timestamp 1681620392
transform 1 0 1196 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1664
timestamp 1681620392
transform 1 0 1180 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1363
timestamp 1681620392
transform 1 0 1188 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1319
timestamp 1681620392
transform 1 0 1228 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1549
timestamp 1681620392
transform 1 0 1236 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1578
timestamp 1681620392
transform 1 0 1236 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1665
timestamp 1681620392
transform 1 0 1196 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1364
timestamp 1681620392
transform 1 0 1212 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_1666
timestamp 1681620392
transform 1 0 1220 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1720
timestamp 1681620392
transform 1 0 1188 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1379
timestamp 1681620392
transform 1 0 1196 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_1721
timestamp 1681620392
transform 1 0 1212 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1380
timestamp 1681620392
transform 1 0 1220 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_1740
timestamp 1681620392
transform 1 0 1188 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_1415
timestamp 1681620392
transform 1 0 1228 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_1579
timestamp 1681620392
transform 1 0 1260 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1667
timestamp 1681620392
transform 1 0 1252 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1288
timestamp 1681620392
transform 1 0 1276 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1289
timestamp 1681620392
transform 1 0 1324 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1320
timestamp 1681620392
transform 1 0 1332 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1580
timestamp 1681620392
transform 1 0 1276 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1581
timestamp 1681620392
transform 1 0 1300 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1582
timestamp 1681620392
transform 1 0 1324 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1583
timestamp 1681620392
transform 1 0 1332 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1722
timestamp 1681620392
transform 1 0 1276 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1381
timestamp 1681620392
transform 1 0 1292 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_1741
timestamp 1681620392
transform 1 0 1268 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_1390
timestamp 1681620392
transform 1 0 1276 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1290
timestamp 1681620392
transform 1 0 1356 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_1550
timestamp 1681620392
transform 1 0 1364 0 1 2145
box -2 -2 2 2
use M3_M2  M3_M2_1321
timestamp 1681620392
transform 1 0 1372 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1584
timestamp 1681620392
transform 1 0 1356 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1585
timestamp 1681620392
transform 1 0 1372 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1668
timestamp 1681620392
transform 1 0 1332 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1669
timestamp 1681620392
transform 1 0 1348 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1723
timestamp 1681620392
transform 1 0 1332 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1391
timestamp 1681620392
transform 1 0 1316 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1392
timestamp 1681620392
transform 1 0 1332 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1291
timestamp 1681620392
transform 1 0 1404 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1292
timestamp 1681620392
transform 1 0 1428 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1293
timestamp 1681620392
transform 1 0 1468 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1322
timestamp 1681620392
transform 1 0 1452 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1323
timestamp 1681620392
transform 1 0 1492 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1586
timestamp 1681620392
transform 1 0 1404 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1587
timestamp 1681620392
transform 1 0 1492 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1670
timestamp 1681620392
transform 1 0 1388 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1365
timestamp 1681620392
transform 1 0 1404 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_1671
timestamp 1681620392
transform 1 0 1452 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1672
timestamp 1681620392
transform 1 0 1484 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1382
timestamp 1681620392
transform 1 0 1388 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1270
timestamp 1681620392
transform 1 0 1516 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_1588
timestamp 1681620392
transform 1 0 1516 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1673
timestamp 1681620392
transform 1 0 1508 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1724
timestamp 1681620392
transform 1 0 1492 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1393
timestamp 1681620392
transform 1 0 1500 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1271
timestamp 1681620392
transform 1 0 1532 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1394
timestamp 1681620392
transform 1 0 1524 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1294
timestamp 1681620392
transform 1 0 1540 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_1589
timestamp 1681620392
transform 1 0 1540 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_1348
timestamp 1681620392
transform 1 0 1612 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_1674
timestamp 1681620392
transform 1 0 1588 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1295
timestamp 1681620392
transform 1 0 1636 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1349
timestamp 1681620392
transform 1 0 1636 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_1675
timestamp 1681620392
transform 1 0 1636 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1590
timestamp 1681620392
transform 1 0 1660 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_1272
timestamp 1681620392
transform 1 0 1668 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_1676
timestamp 1681620392
transform 1 0 1684 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1725
timestamp 1681620392
transform 1 0 1668 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1296
timestamp 1681620392
transform 1 0 1700 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1297
timestamp 1681620392
transform 1 0 1716 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_1591
timestamp 1681620392
transform 1 0 1716 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_1273
timestamp 1681620392
transform 1 0 1732 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1298
timestamp 1681620392
transform 1 0 1796 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1324
timestamp 1681620392
transform 1 0 1796 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1325
timestamp 1681620392
transform 1 0 1812 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1592
timestamp 1681620392
transform 1 0 1732 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_1350
timestamp 1681620392
transform 1 0 1740 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_1593
timestamp 1681620392
transform 1 0 1748 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_1351
timestamp 1681620392
transform 1 0 1764 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_1594
timestamp 1681620392
transform 1 0 1772 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1595
timestamp 1681620392
transform 1 0 1788 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1596
timestamp 1681620392
transform 1 0 1796 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1677
timestamp 1681620392
transform 1 0 1740 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1678
timestamp 1681620392
transform 1 0 1764 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1726
timestamp 1681620392
transform 1 0 1748 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1679
timestamp 1681620392
transform 1 0 1796 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1274
timestamp 1681620392
transform 1 0 1860 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1275
timestamp 1681620392
transform 1 0 1892 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1276
timestamp 1681620392
transform 1 0 1908 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1299
timestamp 1681620392
transform 1 0 1852 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_1597
timestamp 1681620392
transform 1 0 1820 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1598
timestamp 1681620392
transform 1 0 1828 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_1395
timestamp 1681620392
transform 1 0 1804 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1326
timestamp 1681620392
transform 1 0 1908 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1277
timestamp 1681620392
transform 1 0 1956 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1300
timestamp 1681620392
transform 1 0 1964 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_1599
timestamp 1681620392
transform 1 0 1860 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_1352
timestamp 1681620392
transform 1 0 1940 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_1600
timestamp 1681620392
transform 1 0 1948 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_1327
timestamp 1681620392
transform 1 0 1972 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1601
timestamp 1681620392
transform 1 0 1972 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1602
timestamp 1681620392
transform 1 0 1980 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1680
timestamp 1681620392
transform 1 0 1908 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1681
timestamp 1681620392
transform 1 0 1948 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1682
timestamp 1681620392
transform 1 0 1956 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1727
timestamp 1681620392
transform 1 0 1844 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1396
timestamp 1681620392
transform 1 0 1844 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1410
timestamp 1681620392
transform 1 0 1836 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1397
timestamp 1681620392
transform 1 0 1948 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1301
timestamp 1681620392
transform 1 0 2036 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_1603
timestamp 1681620392
transform 1 0 2020 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1604
timestamp 1681620392
transform 1 0 2036 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1683
timestamp 1681620392
transform 1 0 2012 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1728
timestamp 1681620392
transform 1 0 2004 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1398
timestamp 1681620392
transform 1 0 1980 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1411
timestamp 1681620392
transform 1 0 2004 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1353
timestamp 1681620392
transform 1 0 2060 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_1605
timestamp 1681620392
transform 1 0 2140 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1684
timestamp 1681620392
transform 1 0 2084 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1685
timestamp 1681620392
transform 1 0 2124 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1686
timestamp 1681620392
transform 1 0 2132 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1729
timestamp 1681620392
transform 1 0 2124 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1416
timestamp 1681620392
transform 1 0 2092 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1417
timestamp 1681620392
transform 1 0 2132 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_1606
timestamp 1681620392
transform 1 0 2172 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1687
timestamp 1681620392
transform 1 0 2180 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1328
timestamp 1681620392
transform 1 0 2212 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1607
timestamp 1681620392
transform 1 0 2212 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1730
timestamp 1681620392
transform 1 0 2204 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1302
timestamp 1681620392
transform 1 0 2236 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1329
timestamp 1681620392
transform 1 0 2260 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1330
timestamp 1681620392
transform 1 0 2324 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1608
timestamp 1681620392
transform 1 0 2236 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1609
timestamp 1681620392
transform 1 0 2324 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1688
timestamp 1681620392
transform 1 0 2260 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1689
timestamp 1681620392
transform 1 0 2316 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1690
timestamp 1681620392
transform 1 0 2324 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1303
timestamp 1681620392
transform 1 0 2356 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1304
timestamp 1681620392
transform 1 0 2372 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1331
timestamp 1681620392
transform 1 0 2388 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1610
timestamp 1681620392
transform 1 0 2380 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1731
timestamp 1681620392
transform 1 0 2388 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1399
timestamp 1681620392
transform 1 0 2388 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_1732
timestamp 1681620392
transform 1 0 2412 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1400
timestamp 1681620392
transform 1 0 2412 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_1611
timestamp 1681620392
transform 1 0 2436 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_1332
timestamp 1681620392
transform 1 0 2460 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1612
timestamp 1681620392
transform 1 0 2452 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1613
timestamp 1681620392
transform 1 0 2460 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_1278
timestamp 1681620392
transform 1 0 2524 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1279
timestamp 1681620392
transform 1 0 2548 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1333
timestamp 1681620392
transform 1 0 2516 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1614
timestamp 1681620392
transform 1 0 2484 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1615
timestamp 1681620392
transform 1 0 2492 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1616
timestamp 1681620392
transform 1 0 2516 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1691
timestamp 1681620392
transform 1 0 2460 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1692
timestamp 1681620392
transform 1 0 2468 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1693
timestamp 1681620392
transform 1 0 2516 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1733
timestamp 1681620392
transform 1 0 2508 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1401
timestamp 1681620392
transform 1 0 2508 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1305
timestamp 1681620392
transform 1 0 2556 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1306
timestamp 1681620392
transform 1 0 2596 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1334
timestamp 1681620392
transform 1 0 2540 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1335
timestamp 1681620392
transform 1 0 2580 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1307
timestamp 1681620392
transform 1 0 2708 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1336
timestamp 1681620392
transform 1 0 2660 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1337
timestamp 1681620392
transform 1 0 2684 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1617
timestamp 1681620392
transform 1 0 2540 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1618
timestamp 1681620392
transform 1 0 2556 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1619
timestamp 1681620392
transform 1 0 2644 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1694
timestamp 1681620392
transform 1 0 2580 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1366
timestamp 1681620392
transform 1 0 2620 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1354
timestamp 1681620392
transform 1 0 2652 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_1620
timestamp 1681620392
transform 1 0 2660 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1621
timestamp 1681620392
transform 1 0 2676 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1622
timestamp 1681620392
transform 1 0 2684 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1695
timestamp 1681620392
transform 1 0 2636 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1696
timestamp 1681620392
transform 1 0 2652 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1734
timestamp 1681620392
transform 1 0 2540 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1402
timestamp 1681620392
transform 1 0 2628 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1367
timestamp 1681620392
transform 1 0 2660 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1355
timestamp 1681620392
transform 1 0 2700 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1308
timestamp 1681620392
transform 1 0 2732 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_1623
timestamp 1681620392
transform 1 0 2708 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1624
timestamp 1681620392
transform 1 0 2716 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1697
timestamp 1681620392
transform 1 0 2668 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1698
timestamp 1681620392
transform 1 0 2684 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1699
timestamp 1681620392
transform 1 0 2700 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1700
timestamp 1681620392
transform 1 0 2716 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1701
timestamp 1681620392
transform 1 0 2724 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1418
timestamp 1681620392
transform 1 0 2700 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1338
timestamp 1681620392
transform 1 0 2740 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1625
timestamp 1681620392
transform 1 0 2740 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_1403
timestamp 1681620392
transform 1 0 2732 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1309
timestamp 1681620392
transform 1 0 2788 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1339
timestamp 1681620392
transform 1 0 2828 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1626
timestamp 1681620392
transform 1 0 2780 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1627
timestamp 1681620392
transform 1 0 2788 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1628
timestamp 1681620392
transform 1 0 2804 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1702
timestamp 1681620392
transform 1 0 2756 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1703
timestamp 1681620392
transform 1 0 2764 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1383
timestamp 1681620392
transform 1 0 2764 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1368
timestamp 1681620392
transform 1 0 2804 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_1704
timestamp 1681620392
transform 1 0 2820 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_1384
timestamp 1681620392
transform 1 0 2796 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_1735
timestamp 1681620392
transform 1 0 2804 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1412
timestamp 1681620392
transform 1 0 2804 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1419
timestamp 1681620392
transform 1 0 2820 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1280
timestamp 1681620392
transform 1 0 2860 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1281
timestamp 1681620392
transform 1 0 2916 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1340
timestamp 1681620392
transform 1 0 2876 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1341
timestamp 1681620392
transform 1 0 2892 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1342
timestamp 1681620392
transform 1 0 2932 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_1629
timestamp 1681620392
transform 1 0 2844 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1630
timestamp 1681620392
transform 1 0 2860 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1631
timestamp 1681620392
transform 1 0 2868 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_1369
timestamp 1681620392
transform 1 0 2852 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1370
timestamp 1681620392
transform 1 0 2868 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_1632
timestamp 1681620392
transform 1 0 2892 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1633
timestamp 1681620392
transform 1 0 2908 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1705
timestamp 1681620392
transform 1 0 2876 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1736
timestamp 1681620392
transform 1 0 2844 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1282
timestamp 1681620392
transform 1 0 3012 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_1634
timestamp 1681620392
transform 1 0 3012 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1706
timestamp 1681620392
transform 1 0 2932 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1707
timestamp 1681620392
transform 1 0 2996 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1708
timestamp 1681620392
transform 1 0 3004 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1737
timestamp 1681620392
transform 1 0 2892 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1404
timestamp 1681620392
transform 1 0 2892 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_1738
timestamp 1681620392
transform 1 0 2996 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_1413
timestamp 1681620392
transform 1 0 2940 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1405
timestamp 1681620392
transform 1 0 3004 0 1 2105
box -3 -3 3 3
use Project_Top_VIA0  Project_Top_VIA0_18
timestamp 1681620392
transform 1 0 24 0 1 2070
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_93
timestamp 1681620392
transform 1 0 72 0 -1 2170
box -8 -3 104 105
use NAND2X1  NAND2X1_73
timestamp 1681620392
transform 1 0 168 0 -1 2170
box -8 -3 32 105
use AOI22X1  AOI22X1_19
timestamp 1681620392
transform 1 0 192 0 -1 2170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_94
timestamp 1681620392
transform -1 0 328 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_95
timestamp 1681620392
transform 1 0 328 0 -1 2170
box -8 -3 104 105
use OAI21X1  OAI21X1_95
timestamp 1681620392
transform -1 0 456 0 -1 2170
box -8 -3 34 105
use INVX2  INVX2_87
timestamp 1681620392
transform -1 0 472 0 -1 2170
box -9 -3 26 105
use FILL  FILL_304
timestamp 1681620392
transform 1 0 472 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_96
timestamp 1681620392
transform -1 0 576 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_97
timestamp 1681620392
transform 1 0 576 0 -1 2170
box -8 -3 104 105
use OAI21X1  OAI21X1_96
timestamp 1681620392
transform 1 0 672 0 -1 2170
box -8 -3 34 105
use FILL  FILL_307
timestamp 1681620392
transform 1 0 704 0 -1 2170
box -8 -3 16 105
use FILL  FILL_308
timestamp 1681620392
transform 1 0 712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_309
timestamp 1681620392
transform 1 0 720 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_90
timestamp 1681620392
transform -1 0 744 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_91
timestamp 1681620392
transform 1 0 744 0 -1 2170
box -9 -3 26 105
use OAI21X1  OAI21X1_97
timestamp 1681620392
transform 1 0 760 0 -1 2170
box -8 -3 34 105
use FILL  FILL_310
timestamp 1681620392
transform 1 0 792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_311
timestamp 1681620392
transform 1 0 800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_312
timestamp 1681620392
transform 1 0 808 0 -1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_26
timestamp 1681620392
transform 1 0 816 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_76
timestamp 1681620392
transform -1 0 864 0 -1 2170
box -8 -3 32 105
use M3_M2  M3_M2_1420
timestamp 1681620392
transform 1 0 876 0 1 2075
box -3 -3 3 3
use INVX2  INVX2_92
timestamp 1681620392
transform -1 0 880 0 -1 2170
box -9 -3 26 105
use NAND2X1  NAND2X1_77
timestamp 1681620392
transform 1 0 880 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_78
timestamp 1681620392
transform 1 0 904 0 -1 2170
box -8 -3 32 105
use FILL  FILL_314
timestamp 1681620392
transform 1 0 928 0 -1 2170
box -8 -3 16 105
use FILL  FILL_315
timestamp 1681620392
transform 1 0 936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_316
timestamp 1681620392
transform 1 0 944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_325
timestamp 1681620392
transform 1 0 952 0 -1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_92
timestamp 1681620392
transform 1 0 960 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_93
timestamp 1681620392
transform 1 0 984 0 -1 2170
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_102
timestamp 1681620392
transform 1 0 1008 0 -1 2170
box -8 -3 104 105
use NAND3X1  NAND3X1_38
timestamp 1681620392
transform 1 0 1104 0 -1 2170
box -8 -3 40 105
use INVX2  INVX2_97
timestamp 1681620392
transform -1 0 1152 0 -1 2170
box -9 -3 26 105
use FILL  FILL_326
timestamp 1681620392
transform 1 0 1152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_327
timestamp 1681620392
transform 1 0 1160 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_98
timestamp 1681620392
transform 1 0 1168 0 -1 2170
box -9 -3 26 105
use NAND3X1  NAND3X1_39
timestamp 1681620392
transform 1 0 1184 0 -1 2170
box -8 -3 40 105
use INVX2  INVX2_99
timestamp 1681620392
transform -1 0 1232 0 -1 2170
box -9 -3 26 105
use NOR2X1  NOR2X1_28
timestamp 1681620392
transform 1 0 1232 0 -1 2170
box -8 -3 32 105
use M3_M2  M3_M2_1421
timestamp 1681620392
transform 1 0 1268 0 1 2075
box -3 -3 3 3
use FILL  FILL_328
timestamp 1681620392
transform 1 0 1256 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_1422
timestamp 1681620392
transform 1 0 1292 0 1 2075
box -3 -3 3 3
use NAND3X1  NAND3X1_40
timestamp 1681620392
transform 1 0 1264 0 -1 2170
box -8 -3 40 105
use OAI21X1  OAI21X1_106
timestamp 1681620392
transform -1 0 1328 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_107
timestamp 1681620392
transform -1 0 1360 0 -1 2170
box -8 -3 34 105
use OR2X2  OR2X2_0
timestamp 1681620392
transform 1 0 1360 0 -1 2170
box -7 -3 35 105
use DFFNEGX1  DFFNEGX1_103
timestamp 1681620392
transform 1 0 1392 0 -1 2170
box -8 -3 104 105
use OAI21X1  OAI21X1_108
timestamp 1681620392
transform -1 0 1520 0 -1 2170
box -8 -3 34 105
use FILL  FILL_329
timestamp 1681620392
transform 1 0 1520 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_104
timestamp 1681620392
transform 1 0 1528 0 -1 2170
box -8 -3 104 105
use INVX2  INVX2_100
timestamp 1681620392
transform 1 0 1624 0 -1 2170
box -9 -3 26 105
use FILL  FILL_330
timestamp 1681620392
transform 1 0 1640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_331
timestamp 1681620392
transform 1 0 1648 0 -1 2170
box -8 -3 16 105
use FILL  FILL_332
timestamp 1681620392
transform 1 0 1656 0 -1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_109
timestamp 1681620392
transform -1 0 1696 0 -1 2170
box -8 -3 34 105
use FILL  FILL_333
timestamp 1681620392
transform 1 0 1696 0 -1 2170
box -8 -3 16 105
use FILL  FILL_334
timestamp 1681620392
transform 1 0 1704 0 -1 2170
box -8 -3 16 105
use FILL  FILL_335
timestamp 1681620392
transform 1 0 1712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_336
timestamp 1681620392
transform 1 0 1720 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_101
timestamp 1681620392
transform 1 0 1728 0 -1 2170
box -9 -3 26 105
use OAI21X1  OAI21X1_110
timestamp 1681620392
transform -1 0 1776 0 -1 2170
box -8 -3 34 105
use INVX2  INVX2_102
timestamp 1681620392
transform -1 0 1792 0 -1 2170
box -9 -3 26 105
use OAI21X1  OAI21X1_111
timestamp 1681620392
transform 1 0 1792 0 -1 2170
box -8 -3 34 105
use NAND2X1  NAND2X1_94
timestamp 1681620392
transform 1 0 1824 0 -1 2170
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_105
timestamp 1681620392
transform 1 0 1848 0 -1 2170
box -8 -3 104 105
use OAI21X1  OAI21X1_112
timestamp 1681620392
transform 1 0 1944 0 -1 2170
box -8 -3 34 105
use NAND2X1  NAND2X1_95
timestamp 1681620392
transform 1 0 1976 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_96
timestamp 1681620392
transform -1 0 2024 0 -1 2170
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_106
timestamp 1681620392
transform 1 0 2024 0 -1 2170
box -8 -3 104 105
use NAND2X1  NAND2X1_97
timestamp 1681620392
transform -1 0 2144 0 -1 2170
box -8 -3 32 105
use FILL  FILL_337
timestamp 1681620392
transform 1 0 2144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_338
timestamp 1681620392
transform 1 0 2152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_339
timestamp 1681620392
transform 1 0 2160 0 -1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_113
timestamp 1681620392
transform 1 0 2168 0 -1 2170
box -8 -3 34 105
use FILL  FILL_340
timestamp 1681620392
transform 1 0 2200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_354
timestamp 1681620392
transform 1 0 2208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_355
timestamp 1681620392
transform 1 0 2216 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_111
timestamp 1681620392
transform 1 0 2224 0 -1 2170
box -8 -3 104 105
use OAI21X1  OAI21X1_118
timestamp 1681620392
transform 1 0 2320 0 -1 2170
box -8 -3 34 105
use FILL  FILL_356
timestamp 1681620392
transform 1 0 2352 0 -1 2170
box -8 -3 16 105
use FILL  FILL_357
timestamp 1681620392
transform 1 0 2360 0 -1 2170
box -8 -3 16 105
use FILL  FILL_358
timestamp 1681620392
transform 1 0 2368 0 -1 2170
box -8 -3 16 105
use FILL  FILL_359
timestamp 1681620392
transform 1 0 2376 0 -1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_105
timestamp 1681620392
transform -1 0 2408 0 -1 2170
box -8 -3 32 105
use FILL  FILL_360
timestamp 1681620392
transform 1 0 2408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_361
timestamp 1681620392
transform 1 0 2416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_362
timestamp 1681620392
transform 1 0 2424 0 -1 2170
box -8 -3 16 105
use NAND2X1  NAND2X1_106
timestamp 1681620392
transform -1 0 2456 0 -1 2170
box -8 -3 32 105
use OAI21X1  OAI21X1_119
timestamp 1681620392
transform 1 0 2456 0 -1 2170
box -8 -3 34 105
use NAND2X1  NAND2X1_107
timestamp 1681620392
transform 1 0 2488 0 -1 2170
box -8 -3 32 105
use OAI21X1  OAI21X1_120
timestamp 1681620392
transform 1 0 2512 0 -1 2170
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_112
timestamp 1681620392
transform 1 0 2544 0 -1 2170
box -8 -3 104 105
use OAI22X1  OAI22X1_7
timestamp 1681620392
transform 1 0 2640 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_20
timestamp 1681620392
transform -1 0 2720 0 -1 2170
box -8 -3 46 105
use INVX2  INVX2_103
timestamp 1681620392
transform 1 0 2720 0 -1 2170
box -9 -3 26 105
use FILL  FILL_363
timestamp 1681620392
transform 1 0 2736 0 -1 2170
box -8 -3 16 105
use FILL  FILL_364
timestamp 1681620392
transform 1 0 2744 0 -1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_121
timestamp 1681620392
transform 1 0 2752 0 -1 2170
box -8 -3 34 105
use NAND2X1  NAND2X1_108
timestamp 1681620392
transform 1 0 2784 0 -1 2170
box -8 -3 32 105
use OAI21X1  OAI21X1_122
timestamp 1681620392
transform 1 0 2808 0 -1 2170
box -8 -3 34 105
use NAND2X1  NAND2X1_109
timestamp 1681620392
transform -1 0 2864 0 -1 2170
box -8 -3 32 105
use OAI21X1  OAI21X1_123
timestamp 1681620392
transform 1 0 2864 0 -1 2170
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_113
timestamp 1681620392
transform 1 0 2896 0 -1 2170
box -8 -3 104 105
use NAND2X1  NAND2X1_110
timestamp 1681620392
transform -1 0 3016 0 -1 2170
box -8 -3 32 105
use Project_Top_VIA0  Project_Top_VIA0_19
timestamp 1681620392
transform 1 0 3067 0 1 2070
box -10 -3 10 3
use M3_M2  M3_M2_1445
timestamp 1681620392
transform 1 0 68 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1742
timestamp 1681620392
transform 1 0 116 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1755
timestamp 1681620392
transform 1 0 68 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1478
timestamp 1681620392
transform 1 0 84 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_1756
timestamp 1681620392
transform 1 0 92 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1757
timestamp 1681620392
transform 1 0 108 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1446
timestamp 1681620392
transform 1 0 148 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1758
timestamp 1681620392
transform 1 0 132 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1759
timestamp 1681620392
transform 1 0 148 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1760
timestamp 1681620392
transform 1 0 156 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1830
timestamp 1681620392
transform 1 0 84 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1831
timestamp 1681620392
transform 1 0 100 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1832
timestamp 1681620392
transform 1 0 116 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1833
timestamp 1681620392
transform 1 0 164 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1513
timestamp 1681620392
transform 1 0 156 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1546
timestamp 1681620392
transform 1 0 100 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1547
timestamp 1681620392
transform 1 0 116 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1548
timestamp 1681620392
transform 1 0 132 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1423
timestamp 1681620392
transform 1 0 180 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1424
timestamp 1681620392
transform 1 0 196 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1549
timestamp 1681620392
transform 1 0 172 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1447
timestamp 1681620392
transform 1 0 204 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1761
timestamp 1681620392
transform 1 0 196 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1762
timestamp 1681620392
transform 1 0 212 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1834
timestamp 1681620392
transform 1 0 188 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1902
timestamp 1681620392
transform 1 0 220 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_1835
timestamp 1681620392
transform 1 0 244 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1763
timestamp 1681620392
transform 1 0 260 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1764
timestamp 1681620392
transform 1 0 268 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1494
timestamp 1681620392
transform 1 0 260 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_1903
timestamp 1681620392
transform 1 0 260 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_1479
timestamp 1681620392
transform 1 0 292 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_1765
timestamp 1681620392
transform 1 0 316 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1480
timestamp 1681620392
transform 1 0 324 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1448
timestamp 1681620392
transform 1 0 428 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1449
timestamp 1681620392
transform 1 0 476 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1766
timestamp 1681620392
transform 1 0 372 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1495
timestamp 1681620392
transform 1 0 276 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_1836
timestamp 1681620392
transform 1 0 292 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1550
timestamp 1681620392
transform 1 0 268 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1551
timestamp 1681620392
transform 1 0 292 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1481
timestamp 1681620392
transform 1 0 388 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_1767
timestamp 1681620392
transform 1 0 412 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1768
timestamp 1681620392
transform 1 0 468 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1769
timestamp 1681620392
transform 1 0 476 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1837
timestamp 1681620392
transform 1 0 388 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1838
timestamp 1681620392
transform 1 0 484 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1839
timestamp 1681620392
transform 1 0 492 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1450
timestamp 1681620392
transform 1 0 508 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1770
timestamp 1681620392
transform 1 0 508 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1840
timestamp 1681620392
transform 1 0 524 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1451
timestamp 1681620392
transform 1 0 540 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1771
timestamp 1681620392
transform 1 0 540 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1841
timestamp 1681620392
transform 1 0 540 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1842
timestamp 1681620392
transform 1 0 548 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1452
timestamp 1681620392
transform 1 0 564 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1772
timestamp 1681620392
transform 1 0 564 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1453
timestamp 1681620392
transform 1 0 668 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1482
timestamp 1681620392
transform 1 0 588 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_1773
timestamp 1681620392
transform 1 0 636 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1774
timestamp 1681620392
transform 1 0 668 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1775
timestamp 1681620392
transform 1 0 676 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1843
timestamp 1681620392
transform 1 0 588 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1496
timestamp 1681620392
transform 1 0 652 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1454
timestamp 1681620392
transform 1 0 692 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1844
timestamp 1681620392
transform 1 0 684 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1845
timestamp 1681620392
transform 1 0 692 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1776
timestamp 1681620392
transform 1 0 700 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1497
timestamp 1681620392
transform 1 0 700 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_1777
timestamp 1681620392
transform 1 0 748 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1778
timestamp 1681620392
transform 1 0 756 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1846
timestamp 1681620392
transform 1 0 740 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1498
timestamp 1681620392
transform 1 0 756 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1435
timestamp 1681620392
transform 1 0 780 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_1904
timestamp 1681620392
transform 1 0 772 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_1552
timestamp 1681620392
transform 1 0 772 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1436
timestamp 1681620392
transform 1 0 820 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_1779
timestamp 1681620392
transform 1 0 844 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1847
timestamp 1681620392
transform 1 0 836 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1848
timestamp 1681620392
transform 1 0 852 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1514
timestamp 1681620392
transform 1 0 852 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1499
timestamp 1681620392
transform 1 0 876 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_1780
timestamp 1681620392
transform 1 0 900 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1849
timestamp 1681620392
transform 1 0 884 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1850
timestamp 1681620392
transform 1 0 892 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1851
timestamp 1681620392
transform 1 0 900 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1905
timestamp 1681620392
transform 1 0 868 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_1515
timestamp 1681620392
transform 1 0 876 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1516
timestamp 1681620392
transform 1 0 892 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1553
timestamp 1681620392
transform 1 0 884 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_1852
timestamp 1681620392
transform 1 0 924 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1517
timestamp 1681620392
transform 1 0 924 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_1906
timestamp 1681620392
transform 1 0 932 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_1455
timestamp 1681620392
transform 1 0 956 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1781
timestamp 1681620392
transform 1 0 956 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1782
timestamp 1681620392
transform 1 0 964 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1783
timestamp 1681620392
transform 1 0 972 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1853
timestamp 1681620392
transform 1 0 956 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1456
timestamp 1681620392
transform 1 0 1028 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1483
timestamp 1681620392
transform 1 0 1004 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_1784
timestamp 1681620392
transform 1 0 1028 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1785
timestamp 1681620392
transform 1 0 1084 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1854
timestamp 1681620392
transform 1 0 980 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1500
timestamp 1681620392
transform 1 0 988 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_1855
timestamp 1681620392
transform 1 0 1004 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1518
timestamp 1681620392
transform 1 0 980 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_1907
timestamp 1681620392
transform 1 0 988 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_1431
timestamp 1681620392
transform 1 0 1172 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1484
timestamp 1681620392
transform 1 0 1108 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_1786
timestamp 1681620392
transform 1 0 1132 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1787
timestamp 1681620392
transform 1 0 1188 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1788
timestamp 1681620392
transform 1 0 1196 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1856
timestamp 1681620392
transform 1 0 1108 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1519
timestamp 1681620392
transform 1 0 1132 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_1743
timestamp 1681620392
transform 1 0 1236 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1857
timestamp 1681620392
transform 1 0 1244 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1520
timestamp 1681620392
transform 1 0 1244 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_1858
timestamp 1681620392
transform 1 0 1260 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1521
timestamp 1681620392
transform 1 0 1260 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1425
timestamp 1681620392
transform 1 0 1356 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1457
timestamp 1681620392
transform 1 0 1300 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1458
timestamp 1681620392
transform 1 0 1324 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1459
timestamp 1681620392
transform 1 0 1348 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1460
timestamp 1681620392
transform 1 0 1388 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1789
timestamp 1681620392
transform 1 0 1284 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1790
timestamp 1681620392
transform 1 0 1292 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1791
timestamp 1681620392
transform 1 0 1324 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1792
timestamp 1681620392
transform 1 0 1388 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1501
timestamp 1681620392
transform 1 0 1284 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1502
timestamp 1681620392
transform 1 0 1308 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_1859
timestamp 1681620392
transform 1 0 1372 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1437
timestamp 1681620392
transform 1 0 1436 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1461
timestamp 1681620392
transform 1 0 1508 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1744
timestamp 1681620392
transform 1 0 1516 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_1462
timestamp 1681620392
transform 1 0 1532 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1793
timestamp 1681620392
transform 1 0 1460 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1485
timestamp 1681620392
transform 1 0 1492 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_1794
timestamp 1681620392
transform 1 0 1508 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1860
timestamp 1681620392
transform 1 0 1396 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1861
timestamp 1681620392
transform 1 0 1412 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1522
timestamp 1681620392
transform 1 0 1444 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1523
timestamp 1681620392
transform 1 0 1460 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_1795
timestamp 1681620392
transform 1 0 1532 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1862
timestamp 1681620392
transform 1 0 1516 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1524
timestamp 1681620392
transform 1 0 1516 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_1863
timestamp 1681620392
transform 1 0 1540 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1525
timestamp 1681620392
transform 1 0 1540 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_1745
timestamp 1681620392
transform 1 0 1580 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1796
timestamp 1681620392
transform 1 0 1564 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1864
timestamp 1681620392
transform 1 0 1556 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1865
timestamp 1681620392
transform 1 0 1604 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1554
timestamp 1681620392
transform 1 0 1612 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_1797
timestamp 1681620392
transform 1 0 1636 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1463
timestamp 1681620392
transform 1 0 1660 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1427
timestamp 1681620392
transform 1 0 1868 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1464
timestamp 1681620392
transform 1 0 1780 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1465
timestamp 1681620392
transform 1 0 1868 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1798
timestamp 1681620392
transform 1 0 1708 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1799
timestamp 1681620392
transform 1 0 1740 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1800
timestamp 1681620392
transform 1 0 1756 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1801
timestamp 1681620392
transform 1 0 1772 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1486
timestamp 1681620392
transform 1 0 1780 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_1802
timestamp 1681620392
transform 1 0 1788 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1803
timestamp 1681620392
transform 1 0 1820 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1866
timestamp 1681620392
transform 1 0 1644 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1867
timestamp 1681620392
transform 1 0 1660 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1868
timestamp 1681620392
transform 1 0 1748 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1869
timestamp 1681620392
transform 1 0 1764 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1870
timestamp 1681620392
transform 1 0 1780 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1526
timestamp 1681620392
transform 1 0 1644 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1527
timestamp 1681620392
transform 1 0 1708 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1503
timestamp 1681620392
transform 1 0 1788 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1504
timestamp 1681620392
transform 1 0 1820 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_1871
timestamp 1681620392
transform 1 0 1868 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1528
timestamp 1681620392
transform 1 0 1764 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1529
timestamp 1681620392
transform 1 0 1780 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1530
timestamp 1681620392
transform 1 0 1796 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1438
timestamp 1681620392
transform 1 0 1972 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1466
timestamp 1681620392
transform 1 0 1916 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1467
timestamp 1681620392
transform 1 0 1932 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1468
timestamp 1681620392
transform 1 0 1980 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1804
timestamp 1681620392
transform 1 0 1932 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1872
timestamp 1681620392
transform 1 0 1892 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1531
timestamp 1681620392
transform 1 0 1892 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1555
timestamp 1681620392
transform 1 0 1908 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_1805
timestamp 1681620392
transform 1 0 1988 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1873
timestamp 1681620392
transform 1 0 1996 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1746
timestamp 1681620392
transform 1 0 2012 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1806
timestamp 1681620392
transform 1 0 2028 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1556
timestamp 1681620392
transform 1 0 2012 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_1807
timestamp 1681620392
transform 1 0 2044 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1874
timestamp 1681620392
transform 1 0 2036 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1557
timestamp 1681620392
transform 1 0 2036 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_1875
timestamp 1681620392
transform 1 0 2060 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1747
timestamp 1681620392
transform 1 0 2092 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_1487
timestamp 1681620392
transform 1 0 2132 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_1808
timestamp 1681620392
transform 1 0 2156 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1432
timestamp 1681620392
transform 1 0 2252 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1469
timestamp 1681620392
transform 1 0 2260 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1809
timestamp 1681620392
transform 1 0 2204 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1810
timestamp 1681620392
transform 1 0 2268 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1876
timestamp 1681620392
transform 1 0 2092 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1877
timestamp 1681620392
transform 1 0 2108 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1505
timestamp 1681620392
transform 1 0 2156 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1506
timestamp 1681620392
transform 1 0 2188 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1532
timestamp 1681620392
transform 1 0 2108 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_1878
timestamp 1681620392
transform 1 0 2220 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1533
timestamp 1681620392
transform 1 0 2268 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1470
timestamp 1681620392
transform 1 0 2356 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1471
timestamp 1681620392
transform 1 0 2436 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1748
timestamp 1681620392
transform 1 0 2460 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1811
timestamp 1681620392
transform 1 0 2324 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1812
timestamp 1681620392
transform 1 0 2332 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1488
timestamp 1681620392
transform 1 0 2340 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_1813
timestamp 1681620392
transform 1 0 2348 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1507
timestamp 1681620392
transform 1 0 2324 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_1814
timestamp 1681620392
transform 1 0 2420 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1815
timestamp 1681620392
transform 1 0 2452 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1472
timestamp 1681620392
transform 1 0 2476 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1816
timestamp 1681620392
transform 1 0 2476 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1879
timestamp 1681620392
transform 1 0 2340 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1880
timestamp 1681620392
transform 1 0 2356 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1881
timestamp 1681620392
transform 1 0 2372 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1882
timestamp 1681620392
transform 1 0 2460 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1534
timestamp 1681620392
transform 1 0 2340 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1535
timestamp 1681620392
transform 1 0 2420 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1536
timestamp 1681620392
transform 1 0 2460 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1558
timestamp 1681620392
transform 1 0 2444 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_1883
timestamp 1681620392
transform 1 0 2484 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1749
timestamp 1681620392
transform 1 0 2500 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1750
timestamp 1681620392
transform 1 0 2508 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_1489
timestamp 1681620392
transform 1 0 2500 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_1817
timestamp 1681620392
transform 1 0 2508 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1508
timestamp 1681620392
transform 1 0 2500 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1559
timestamp 1681620392
transform 1 0 2492 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1473
timestamp 1681620392
transform 1 0 2540 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1490
timestamp 1681620392
transform 1 0 2532 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_1884
timestamp 1681620392
transform 1 0 2548 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1537
timestamp 1681620392
transform 1 0 2548 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1426
timestamp 1681620392
transform 1 0 2612 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1474
timestamp 1681620392
transform 1 0 2588 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1818
timestamp 1681620392
transform 1 0 2588 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1819
timestamp 1681620392
transform 1 0 2644 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1885
timestamp 1681620392
transform 1 0 2564 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1509
timestamp 1681620392
transform 1 0 2588 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1510
timestamp 1681620392
transform 1 0 2612 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_1886
timestamp 1681620392
transform 1 0 2652 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1538
timestamp 1681620392
transform 1 0 2596 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1539
timestamp 1681620392
transform 1 0 2644 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1439
timestamp 1681620392
transform 1 0 2692 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_1887
timestamp 1681620392
transform 1 0 2684 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1475
timestamp 1681620392
transform 1 0 2708 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1820
timestamp 1681620392
transform 1 0 2708 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1433
timestamp 1681620392
transform 1 0 2748 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1434
timestamp 1681620392
transform 1 0 2764 0 1 2045
box -3 -3 3 3
use M2_M1  M2_M1_1751
timestamp 1681620392
transform 1 0 2748 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1821
timestamp 1681620392
transform 1 0 2732 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1491
timestamp 1681620392
transform 1 0 2740 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_1888
timestamp 1681620392
transform 1 0 2716 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1889
timestamp 1681620392
transform 1 0 2724 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1511
timestamp 1681620392
transform 1 0 2740 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1440
timestamp 1681620392
transform 1 0 2780 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1441
timestamp 1681620392
transform 1 0 2796 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1442
timestamp 1681620392
transform 1 0 2812 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_1752
timestamp 1681620392
transform 1 0 2780 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1822
timestamp 1681620392
transform 1 0 2764 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1492
timestamp 1681620392
transform 1 0 2788 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_1890
timestamp 1681620392
transform 1 0 2748 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1891
timestamp 1681620392
transform 1 0 2756 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1512
timestamp 1681620392
transform 1 0 2764 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_1892
timestamp 1681620392
transform 1 0 2780 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1893
timestamp 1681620392
transform 1 0 2788 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1894
timestamp 1681620392
transform 1 0 2804 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1540
timestamp 1681620392
transform 1 0 2780 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_1908
timestamp 1681620392
transform 1 0 2788 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_1541
timestamp 1681620392
transform 1 0 2796 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1542
timestamp 1681620392
transform 1 0 2812 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1560
timestamp 1681620392
transform 1 0 2756 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1561
timestamp 1681620392
transform 1 0 2788 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_1823
timestamp 1681620392
transform 1 0 2828 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1895
timestamp 1681620392
transform 1 0 2820 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1896
timestamp 1681620392
transform 1 0 2828 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1476
timestamp 1681620392
transform 1 0 2844 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1824
timestamp 1681620392
transform 1 0 2836 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1825
timestamp 1681620392
transform 1 0 2844 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1897
timestamp 1681620392
transform 1 0 2844 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1543
timestamp 1681620392
transform 1 0 2844 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1428
timestamp 1681620392
transform 1 0 2884 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1429
timestamp 1681620392
transform 1 0 2908 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1430
timestamp 1681620392
transform 1 0 2932 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1443
timestamp 1681620392
transform 1 0 2868 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1444
timestamp 1681620392
transform 1 0 2972 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_1753
timestamp 1681620392
transform 1 0 2868 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_1477
timestamp 1681620392
transform 1 0 2908 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_1754
timestamp 1681620392
transform 1 0 2988 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1826
timestamp 1681620392
transform 1 0 2916 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1827
timestamp 1681620392
transform 1 0 2964 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1828
timestamp 1681620392
transform 1 0 2972 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_1493
timestamp 1681620392
transform 1 0 2980 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_1829
timestamp 1681620392
transform 1 0 2996 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1898
timestamp 1681620392
transform 1 0 2868 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1899
timestamp 1681620392
transform 1 0 2884 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1900
timestamp 1681620392
transform 1 0 2972 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_1544
timestamp 1681620392
transform 1 0 2868 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1545
timestamp 1681620392
transform 1 0 2916 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_1901
timestamp 1681620392
transform 1 0 3012 0 1 2005
box -2 -2 2 2
use Project_Top_VIA0  Project_Top_VIA0_20
timestamp 1681620392
transform 1 0 48 0 1 1970
box -10 -3 10 3
use AOI22X1  AOI22X1_21
timestamp 1681620392
transform 1 0 72 0 1 1970
box -8 -3 46 105
use OAI21X1  OAI21X1_124
timestamp 1681620392
transform -1 0 144 0 1 1970
box -8 -3 34 105
use INVX2  INVX2_104
timestamp 1681620392
transform -1 0 160 0 1 1970
box -9 -3 26 105
use FILL  FILL_365
timestamp 1681620392
transform 1 0 160 0 1 1970
box -8 -3 16 105
use FILL  FILL_366
timestamp 1681620392
transform 1 0 168 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_1562
timestamp 1681620392
transform 1 0 188 0 1 1975
box -3 -3 3 3
use AOI22X1  AOI22X1_22
timestamp 1681620392
transform -1 0 216 0 1 1970
box -8 -3 46 105
use M3_M2  M3_M2_1563
timestamp 1681620392
transform 1 0 236 0 1 1975
box -3 -3 3 3
use NOR2X1  NOR2X1_30
timestamp 1681620392
transform 1 0 216 0 1 1970
box -8 -3 32 105
use FILL  FILL_373
timestamp 1681620392
transform 1 0 240 0 1 1970
box -8 -3 16 105
use FILL  FILL_375
timestamp 1681620392
transform 1 0 248 0 1 1970
box -8 -3 16 105
use FILL  FILL_377
timestamp 1681620392
transform 1 0 256 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_106
timestamp 1681620392
transform 1 0 264 0 1 1970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_114
timestamp 1681620392
transform 1 0 280 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_115
timestamp 1681620392
transform 1 0 376 0 1 1970
box -8 -3 104 105
use INVX2  INVX2_107
timestamp 1681620392
transform -1 0 488 0 1 1970
box -9 -3 26 105
use FILL  FILL_379
timestamp 1681620392
transform 1 0 488 0 1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_125
timestamp 1681620392
transform 1 0 496 0 1 1970
box -8 -3 34 105
use INVX2  INVX2_108
timestamp 1681620392
transform -1 0 544 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_109
timestamp 1681620392
transform 1 0 544 0 1 1970
box -9 -3 26 105
use FILL  FILL_380
timestamp 1681620392
transform 1 0 560 0 1 1970
box -8 -3 16 105
use FILL  FILL_381
timestamp 1681620392
transform 1 0 568 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_1564
timestamp 1681620392
transform 1 0 660 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1565
timestamp 1681620392
transform 1 0 676 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_116
timestamp 1681620392
transform 1 0 576 0 1 1970
box -8 -3 104 105
use INVX2  INVX2_110
timestamp 1681620392
transform -1 0 688 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_111
timestamp 1681620392
transform 1 0 688 0 1 1970
box -9 -3 26 105
use FILL  FILL_382
timestamp 1681620392
transform 1 0 704 0 1 1970
box -8 -3 16 105
use FILL  FILL_383
timestamp 1681620392
transform 1 0 712 0 1 1970
box -8 -3 16 105
use FILL  FILL_384
timestamp 1681620392
transform 1 0 720 0 1 1970
box -8 -3 16 105
use FILL  FILL_385
timestamp 1681620392
transform 1 0 728 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_112
timestamp 1681620392
transform 1 0 736 0 1 1970
box -9 -3 26 105
use NOR2X1  NOR2X1_32
timestamp 1681620392
transform -1 0 776 0 1 1970
box -8 -3 32 105
use FILL  FILL_386
timestamp 1681620392
transform 1 0 776 0 1 1970
box -8 -3 16 105
use FILL  FILL_387
timestamp 1681620392
transform 1 0 784 0 1 1970
box -8 -3 16 105
use FILL  FILL_388
timestamp 1681620392
transform 1 0 792 0 1 1970
box -8 -3 16 105
use FILL  FILL_389
timestamp 1681620392
transform 1 0 800 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_1566
timestamp 1681620392
transform 1 0 820 0 1 1975
box -3 -3 3 3
use FILL  FILL_390
timestamp 1681620392
transform 1 0 808 0 1 1970
box -8 -3 16 105
use FILL  FILL_391
timestamp 1681620392
transform 1 0 816 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_25
timestamp 1681620392
transform 1 0 824 0 1 1970
box -8 -3 46 105
use FILL  FILL_392
timestamp 1681620392
transform 1 0 864 0 1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_33
timestamp 1681620392
transform 1 0 872 0 1 1970
box -8 -3 32 105
use AOI21X1  AOI21X1_8
timestamp 1681620392
transform 1 0 896 0 1 1970
box -7 -3 39 105
use FILL  FILL_393
timestamp 1681620392
transform 1 0 928 0 1 1970
box -8 -3 16 105
use FILL  FILL_394
timestamp 1681620392
transform 1 0 936 0 1 1970
box -8 -3 16 105
use FILL  FILL_395
timestamp 1681620392
transform 1 0 944 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_113
timestamp 1681620392
transform 1 0 952 0 1 1970
box -9 -3 26 105
use NOR2X1  NOR2X1_34
timestamp 1681620392
transform -1 0 992 0 1 1970
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_117
timestamp 1681620392
transform 1 0 992 0 1 1970
box -8 -3 104 105
use FILL  FILL_396
timestamp 1681620392
transform 1 0 1088 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_118
timestamp 1681620392
transform 1 0 1096 0 1 1970
box -8 -3 104 105
use BUFX2  BUFX2_13
timestamp 1681620392
transform 1 0 1192 0 1 1970
box -5 -3 28 105
use FILL  FILL_397
timestamp 1681620392
transform 1 0 1216 0 1 1970
box -8 -3 16 105
use FILL  FILL_398
timestamp 1681620392
transform 1 0 1224 0 1 1970
box -8 -3 16 105
use FILL  FILL_399
timestamp 1681620392
transform 1 0 1232 0 1 1970
box -8 -3 16 105
use NAND2X1  NAND2X1_111
timestamp 1681620392
transform -1 0 1264 0 1 1970
box -8 -3 32 105
use FILL  FILL_400
timestamp 1681620392
transform 1 0 1264 0 1 1970
box -8 -3 16 105
use FILL  FILL_401
timestamp 1681620392
transform 1 0 1272 0 1 1970
box -8 -3 16 105
use FILL  FILL_402
timestamp 1681620392
transform 1 0 1280 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_119
timestamp 1681620392
transform -1 0 1384 0 1 1970
box -8 -3 104 105
use INVX2  INVX2_114
timestamp 1681620392
transform -1 0 1400 0 1 1970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_120
timestamp 1681620392
transform 1 0 1400 0 1 1970
box -8 -3 104 105
use INVX2  INVX2_115
timestamp 1681620392
transform 1 0 1496 0 1 1970
box -9 -3 26 105
use OAI21X1  OAI21X1_126
timestamp 1681620392
transform -1 0 1544 0 1 1970
box -8 -3 34 105
use FILL  FILL_403
timestamp 1681620392
transform 1 0 1544 0 1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_130
timestamp 1681620392
transform 1 0 1552 0 1 1970
box -8 -3 34 105
use INVX2  INVX2_125
timestamp 1681620392
transform 1 0 1584 0 1 1970
box -9 -3 26 105
use FILL  FILL_421
timestamp 1681620392
transform 1 0 1600 0 1 1970
box -8 -3 16 105
use FILL  FILL_425
timestamp 1681620392
transform 1 0 1608 0 1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_132
timestamp 1681620392
transform -1 0 1648 0 1 1970
box -8 -3 34 105
use M3_M2  M3_M2_1567
timestamp 1681620392
transform 1 0 1660 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_124
timestamp 1681620392
transform 1 0 1648 0 1 1970
box -8 -3 104 105
use M3_M2  M3_M2_1568
timestamp 1681620392
transform 1 0 1772 0 1 1975
box -3 -3 3 3
use OAI22X1  OAI22X1_12
timestamp 1681620392
transform 1 0 1744 0 1 1970
box -8 -3 46 105
use M3_M2  M3_M2_1569
timestamp 1681620392
transform 1 0 1796 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1570
timestamp 1681620392
transform 1 0 1836 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1571
timestamp 1681620392
transform 1 0 1868 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_125
timestamp 1681620392
transform -1 0 1880 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_126
timestamp 1681620392
transform 1 0 1880 0 1 1970
box -8 -3 104 105
use INVX2  INVX2_126
timestamp 1681620392
transform 1 0 1976 0 1 1970
box -9 -3 26 105
use FILL  FILL_426
timestamp 1681620392
transform 1 0 1992 0 1 1970
box -8 -3 16 105
use FILL  FILL_427
timestamp 1681620392
transform 1 0 2000 0 1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_133
timestamp 1681620392
transform -1 0 2040 0 1 1970
box -8 -3 34 105
use FILL  FILL_428
timestamp 1681620392
transform 1 0 2040 0 1 1970
box -8 -3 16 105
use FILL  FILL_429
timestamp 1681620392
transform 1 0 2048 0 1 1970
box -8 -3 16 105
use FILL  FILL_430
timestamp 1681620392
transform 1 0 2056 0 1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_134
timestamp 1681620392
transform 1 0 2064 0 1 1970
box -8 -3 34 105
use M3_M2  M3_M2_1572
timestamp 1681620392
transform 1 0 2180 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_127
timestamp 1681620392
transform 1 0 2096 0 1 1970
box -8 -3 104 105
use INVX2  INVX2_127
timestamp 1681620392
transform 1 0 2192 0 1 1970
box -9 -3 26 105
use M3_M2  M3_M2_1573
timestamp 1681620392
transform 1 0 2276 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_128
timestamp 1681620392
transform 1 0 2208 0 1 1970
box -8 -3 104 105
use INVX2  INVX2_128
timestamp 1681620392
transform 1 0 2304 0 1 1970
box -9 -3 26 105
use M3_M2  M3_M2_1574
timestamp 1681620392
transform 1 0 2340 0 1 1975
box -3 -3 3 3
use OAI22X1  OAI22X1_13
timestamp 1681620392
transform 1 0 2320 0 1 1970
box -8 -3 46 105
use M3_M2  M3_M2_1575
timestamp 1681620392
transform 1 0 2372 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1576
timestamp 1681620392
transform 1 0 2388 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1577
timestamp 1681620392
transform 1 0 2404 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_129
timestamp 1681620392
transform 1 0 2360 0 1 1970
box -8 -3 104 105
use OAI21X1  OAI21X1_135
timestamp 1681620392
transform -1 0 2488 0 1 1970
box -8 -3 34 105
use FILL  FILL_431
timestamp 1681620392
transform 1 0 2488 0 1 1970
box -8 -3 16 105
use FILL  FILL_432
timestamp 1681620392
transform 1 0 2496 0 1 1970
box -8 -3 16 105
use NAND2X1  NAND2X1_114
timestamp 1681620392
transform -1 0 2528 0 1 1970
box -8 -3 32 105
use FILL  FILL_433
timestamp 1681620392
transform 1 0 2528 0 1 1970
box -8 -3 16 105
use FILL  FILL_449
timestamp 1681620392
transform 1 0 2536 0 1 1970
box -8 -3 16 105
use FILL  FILL_451
timestamp 1681620392
transform 1 0 2544 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_133
timestamp 1681620392
transform 1 0 2552 0 1 1970
box -8 -3 104 105
use FILL  FILL_452
timestamp 1681620392
transform 1 0 2648 0 1 1970
box -8 -3 16 105
use FILL  FILL_455
timestamp 1681620392
transform 1 0 2656 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_133
timestamp 1681620392
transform 1 0 2664 0 1 1970
box -9 -3 26 105
use OAI21X1  OAI21X1_138
timestamp 1681620392
transform -1 0 2712 0 1 1970
box -8 -3 34 105
use FILL  FILL_457
timestamp 1681620392
transform 1 0 2712 0 1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_139
timestamp 1681620392
transform 1 0 2720 0 1 1970
box -8 -3 34 105
use M3_M2  M3_M2_1578
timestamp 1681620392
transform 1 0 2764 0 1 1975
box -3 -3 3 3
use OAI21X1  OAI21X1_140
timestamp 1681620392
transform 1 0 2752 0 1 1970
box -8 -3 34 105
use NOR2X1  NOR2X1_38
timestamp 1681620392
transform 1 0 2784 0 1 1970
box -8 -3 32 105
use INVX2  INVX2_134
timestamp 1681620392
transform -1 0 2824 0 1 1970
box -9 -3 26 105
use M3_M2  M3_M2_1579
timestamp 1681620392
transform 1 0 2852 0 1 1975
box -3 -3 3 3
use INVX2  INVX2_135
timestamp 1681620392
transform 1 0 2824 0 1 1970
box -9 -3 26 105
use OAI21X1  OAI21X1_141
timestamp 1681620392
transform 1 0 2840 0 1 1970
box -8 -3 34 105
use M3_M2  M3_M2_1580
timestamp 1681620392
transform 1 0 2892 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_135
timestamp 1681620392
transform 1 0 2872 0 1 1970
box -8 -3 104 105
use NAND2X1  NAND2X1_117
timestamp 1681620392
transform 1 0 2968 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_118
timestamp 1681620392
transform -1 0 3016 0 1 1970
box -8 -3 32 105
use Project_Top_VIA0  Project_Top_VIA0_21
timestamp 1681620392
transform 1 0 3043 0 1 1970
box -10 -3 10 3
use M3_M2  M3_M2_1596
timestamp 1681620392
transform 1 0 84 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_1916
timestamp 1681620392
transform 1 0 84 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2004
timestamp 1681620392
transform 1 0 84 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1745
timestamp 1681620392
transform 1 0 84 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1621
timestamp 1681620392
transform 1 0 108 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1597
timestamp 1681620392
transform 1 0 132 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_1917
timestamp 1681620392
transform 1 0 116 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1663
timestamp 1681620392
transform 1 0 124 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1918
timestamp 1681620392
transform 1 0 132 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2005
timestamp 1681620392
transform 1 0 108 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2006
timestamp 1681620392
transform 1 0 124 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2007
timestamp 1681620392
transform 1 0 132 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1713
timestamp 1681620392
transform 1 0 132 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1598
timestamp 1681620392
transform 1 0 188 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_1919
timestamp 1681620392
transform 1 0 172 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1664
timestamp 1681620392
transform 1 0 180 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_2008
timestamp 1681620392
transform 1 0 164 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1622
timestamp 1681620392
transform 1 0 204 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1909
timestamp 1681620392
transform 1 0 220 0 1 1945
box -2 -2 2 2
use M3_M2  M3_M2_1665
timestamp 1681620392
transform 1 0 196 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_2009
timestamp 1681620392
transform 1 0 188 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2010
timestamp 1681620392
transform 1 0 196 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1666
timestamp 1681620392
transform 1 0 220 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1599
timestamp 1681620392
transform 1 0 244 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_1910
timestamp 1681620392
transform 1 0 236 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1920
timestamp 1681620392
transform 1 0 228 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2011
timestamp 1681620392
transform 1 0 220 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1714
timestamp 1681620392
transform 1 0 204 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1765
timestamp 1681620392
transform 1 0 220 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_1921
timestamp 1681620392
transform 1 0 244 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1667
timestamp 1681620392
transform 1 0 252 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1581
timestamp 1681620392
transform 1 0 276 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1668
timestamp 1681620392
transform 1 0 276 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1582
timestamp 1681620392
transform 1 0 316 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1600
timestamp 1681620392
transform 1 0 332 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1623
timestamp 1681620392
transform 1 0 324 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1911
timestamp 1681620392
transform 1 0 332 0 1 1945
box -2 -2 2 2
use M3_M2  M3_M2_1624
timestamp 1681620392
transform 1 0 356 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1922
timestamp 1681620392
transform 1 0 292 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1923
timestamp 1681620392
transform 1 0 308 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1924
timestamp 1681620392
transform 1 0 324 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1925
timestamp 1681620392
transform 1 0 348 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1926
timestamp 1681620392
transform 1 0 356 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2012
timestamp 1681620392
transform 1 0 284 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1687
timestamp 1681620392
transform 1 0 292 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2013
timestamp 1681620392
transform 1 0 300 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2014
timestamp 1681620392
transform 1 0 316 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2015
timestamp 1681620392
transform 1 0 332 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1688
timestamp 1681620392
transform 1 0 348 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2016
timestamp 1681620392
transform 1 0 356 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1715
timestamp 1681620392
transform 1 0 316 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1716
timestamp 1681620392
transform 1 0 332 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1766
timestamp 1681620392
transform 1 0 284 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1775
timestamp 1681620392
transform 1 0 292 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1776
timestamp 1681620392
transform 1 0 340 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1625
timestamp 1681620392
transform 1 0 372 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1626
timestamp 1681620392
transform 1 0 404 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1927
timestamp 1681620392
transform 1 0 412 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2017
timestamp 1681620392
transform 1 0 388 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2092
timestamp 1681620392
transform 1 0 380 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2116
timestamp 1681620392
transform 1 0 380 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_1777
timestamp 1681620392
transform 1 0 380 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1627
timestamp 1681620392
transform 1 0 436 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1912
timestamp 1681620392
transform 1 0 444 0 1 1945
box -2 -2 2 2
use M3_M2  M3_M2_1583
timestamp 1681620392
transform 1 0 556 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1601
timestamp 1681620392
transform 1 0 500 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1602
timestamp 1681620392
transform 1 0 516 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1603
timestamp 1681620392
transform 1 0 548 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1628
timestamp 1681620392
transform 1 0 492 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1928
timestamp 1681620392
transform 1 0 436 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1929
timestamp 1681620392
transform 1 0 452 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2018
timestamp 1681620392
transform 1 0 428 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1669
timestamp 1681620392
transform 1 0 476 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1930
timestamp 1681620392
transform 1 0 500 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1689
timestamp 1681620392
transform 1 0 452 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2019
timestamp 1681620392
transform 1 0 468 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2020
timestamp 1681620392
transform 1 0 484 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1717
timestamp 1681620392
transform 1 0 436 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1746
timestamp 1681620392
transform 1 0 428 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1747
timestamp 1681620392
transform 1 0 444 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_1913
timestamp 1681620392
transform 1 0 564 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1931
timestamp 1681620392
transform 1 0 516 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1932
timestamp 1681620392
transform 1 0 524 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1670
timestamp 1681620392
transform 1 0 532 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1933
timestamp 1681620392
transform 1 0 540 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1934
timestamp 1681620392
transform 1 0 556 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1935
timestamp 1681620392
transform 1 0 564 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2021
timestamp 1681620392
transform 1 0 516 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1690
timestamp 1681620392
transform 1 0 524 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2022
timestamp 1681620392
transform 1 0 532 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2023
timestamp 1681620392
transform 1 0 548 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2093
timestamp 1681620392
transform 1 0 476 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2094
timestamp 1681620392
transform 1 0 492 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_1748
timestamp 1681620392
transform 1 0 476 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1767
timestamp 1681620392
transform 1 0 468 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1718
timestamp 1681620392
transform 1 0 516 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1691
timestamp 1681620392
transform 1 0 564 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1749
timestamp 1681620392
transform 1 0 532 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1750
timestamp 1681620392
transform 1 0 556 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1768
timestamp 1681620392
transform 1 0 548 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1584
timestamp 1681620392
transform 1 0 588 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_1936
timestamp 1681620392
transform 1 0 588 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2024
timestamp 1681620392
transform 1 0 580 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1604
timestamp 1681620392
transform 1 0 620 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1629
timestamp 1681620392
transform 1 0 628 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1937
timestamp 1681620392
transform 1 0 628 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2025
timestamp 1681620392
transform 1 0 612 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1719
timestamp 1681620392
transform 1 0 612 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_2095
timestamp 1681620392
transform 1 0 628 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_1769
timestamp 1681620392
transform 1 0 580 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1605
timestamp 1681620392
transform 1 0 684 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_1914
timestamp 1681620392
transform 1 0 684 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1938
timestamp 1681620392
transform 1 0 636 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1939
timestamp 1681620392
transform 1 0 660 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1940
timestamp 1681620392
transform 1 0 668 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2026
timestamp 1681620392
transform 1 0 652 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1692
timestamp 1681620392
transform 1 0 668 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_1941
timestamp 1681620392
transform 1 0 692 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1942
timestamp 1681620392
transform 1 0 716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2027
timestamp 1681620392
transform 1 0 676 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2028
timestamp 1681620392
transform 1 0 708 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2096
timestamp 1681620392
transform 1 0 636 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_1720
timestamp 1681620392
transform 1 0 644 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1751
timestamp 1681620392
transform 1 0 628 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1721
timestamp 1681620392
transform 1 0 700 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1770
timestamp 1681620392
transform 1 0 692 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1585
timestamp 1681620392
transform 1 0 788 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1630
timestamp 1681620392
transform 1 0 796 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1915
timestamp 1681620392
transform 1 0 836 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1943
timestamp 1681620392
transform 1 0 820 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1671
timestamp 1681620392
transform 1 0 836 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1606
timestamp 1681620392
transform 1 0 852 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1607
timestamp 1681620392
transform 1 0 892 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_1944
timestamp 1681620392
transform 1 0 844 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2029
timestamp 1681620392
transform 1 0 732 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2030
timestamp 1681620392
transform 1 0 740 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2031
timestamp 1681620392
transform 1 0 796 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1672
timestamp 1681620392
transform 1 0 852 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1673
timestamp 1681620392
transform 1 0 884 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_2032
timestamp 1681620392
transform 1 0 860 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2033
timestamp 1681620392
transform 1 0 868 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2034
timestamp 1681620392
transform 1 0 884 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1722
timestamp 1681620392
transform 1 0 860 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_2097
timestamp 1681620392
transform 1 0 876 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_1723
timestamp 1681620392
transform 1 0 884 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_2098
timestamp 1681620392
transform 1 0 900 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2117
timestamp 1681620392
transform 1 0 884 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_1608
timestamp 1681620392
transform 1 0 932 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1609
timestamp 1681620392
transform 1 0 972 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1631
timestamp 1681620392
transform 1 0 948 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1632
timestamp 1681620392
transform 1 0 964 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1945
timestamp 1681620392
transform 1 0 932 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1674
timestamp 1681620392
transform 1 0 940 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1633
timestamp 1681620392
transform 1 0 1012 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1946
timestamp 1681620392
transform 1 0 948 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1947
timestamp 1681620392
transform 1 0 964 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1948
timestamp 1681620392
transform 1 0 972 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1949
timestamp 1681620392
transform 1 0 980 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1950
timestamp 1681620392
transform 1 0 996 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1951
timestamp 1681620392
transform 1 0 1012 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2035
timestamp 1681620392
transform 1 0 940 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2036
timestamp 1681620392
transform 1 0 972 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1724
timestamp 1681620392
transform 1 0 972 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1778
timestamp 1681620392
transform 1 0 956 0 1 1885
box -3 -3 3 3
use M2_M1  M2_M1_2037
timestamp 1681620392
transform 1 0 988 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1771
timestamp 1681620392
transform 1 0 980 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1693
timestamp 1681620392
transform 1 0 1028 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2099
timestamp 1681620392
transform 1 0 1020 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_1752
timestamp 1681620392
transform 1 0 1020 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1779
timestamp 1681620392
transform 1 0 1020 0 1 1885
box -3 -3 3 3
use M2_M1  M2_M1_2038
timestamp 1681620392
transform 1 0 1044 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1675
timestamp 1681620392
transform 1 0 1076 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1952
timestamp 1681620392
transform 1 0 1084 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1694
timestamp 1681620392
transform 1 0 1060 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2039
timestamp 1681620392
transform 1 0 1068 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1725
timestamp 1681620392
transform 1 0 1060 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_2100
timestamp 1681620392
transform 1 0 1076 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2118
timestamp 1681620392
transform 1 0 1060 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_1780
timestamp 1681620392
transform 1 0 1084 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1610
timestamp 1681620392
transform 1 0 1108 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_1953
timestamp 1681620392
transform 1 0 1108 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1676
timestamp 1681620392
transform 1 0 1116 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_2040
timestamp 1681620392
transform 1 0 1108 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2041
timestamp 1681620392
transform 1 0 1116 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2101
timestamp 1681620392
transform 1 0 1124 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_1753
timestamp 1681620392
transform 1 0 1124 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1781
timestamp 1681620392
transform 1 0 1124 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1586
timestamp 1681620392
transform 1 0 1172 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1587
timestamp 1681620392
transform 1 0 1196 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1611
timestamp 1681620392
transform 1 0 1196 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1634
timestamp 1681620392
transform 1 0 1164 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1635
timestamp 1681620392
transform 1 0 1188 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1954
timestamp 1681620392
transform 1 0 1164 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1677
timestamp 1681620392
transform 1 0 1172 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_2042
timestamp 1681620392
transform 1 0 1140 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1695
timestamp 1681620392
transform 1 0 1156 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2043
timestamp 1681620392
transform 1 0 1164 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1696
timestamp 1681620392
transform 1 0 1180 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2044
timestamp 1681620392
transform 1 0 1188 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2102
timestamp 1681620392
transform 1 0 1156 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2103
timestamp 1681620392
transform 1 0 1180 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2119
timestamp 1681620392
transform 1 0 1148 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_1754
timestamp 1681620392
transform 1 0 1180 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_2045
timestamp 1681620392
transform 1 0 1220 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2104
timestamp 1681620392
transform 1 0 1204 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2105
timestamp 1681620392
transform 1 0 1212 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2120
timestamp 1681620392
transform 1 0 1196 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_1782
timestamp 1681620392
transform 1 0 1156 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1783
timestamp 1681620392
transform 1 0 1180 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1726
timestamp 1681620392
transform 1 0 1220 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1588
timestamp 1681620392
transform 1 0 1268 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_1955
timestamp 1681620392
transform 1 0 1356 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2046
timestamp 1681620392
transform 1 0 1260 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2047
timestamp 1681620392
transform 1 0 1276 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2048
timestamp 1681620392
transform 1 0 1308 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2106
timestamp 1681620392
transform 1 0 1236 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2107
timestamp 1681620392
transform 1 0 1244 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_1727
timestamp 1681620392
transform 1 0 1260 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1697
timestamp 1681620392
transform 1 0 1356 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2108
timestamp 1681620392
transform 1 0 1268 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2121
timestamp 1681620392
transform 1 0 1228 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_1755
timestamp 1681620392
transform 1 0 1236 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1772
timestamp 1681620392
transform 1 0 1244 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_2122
timestamp 1681620392
transform 1 0 1268 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_1756
timestamp 1681620392
transform 1 0 1276 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1784
timestamp 1681620392
transform 1 0 1252 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1636
timestamp 1681620392
transform 1 0 1388 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1637
timestamp 1681620392
transform 1 0 1412 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1956
timestamp 1681620392
transform 1 0 1388 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2049
timestamp 1681620392
transform 1 0 1436 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1728
timestamp 1681620392
transform 1 0 1436 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1785
timestamp 1681620392
transform 1 0 1396 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1698
timestamp 1681620392
transform 1 0 1476 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2050
timestamp 1681620392
transform 1 0 1508 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1729
timestamp 1681620392
transform 1 0 1508 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_2051
timestamp 1681620392
transform 1 0 1524 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2109
timestamp 1681620392
transform 1 0 1532 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_1612
timestamp 1681620392
transform 1 0 1564 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1638
timestamp 1681620392
transform 1 0 1556 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_2110
timestamp 1681620392
transform 1 0 1572 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_1639
timestamp 1681620392
transform 1 0 1596 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1957
timestamp 1681620392
transform 1 0 1596 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1699
timestamp 1681620392
transform 1 0 1596 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2052
timestamp 1681620392
transform 1 0 1604 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1786
timestamp 1681620392
transform 1 0 1604 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1640
timestamp 1681620392
transform 1 0 1628 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1958
timestamp 1681620392
transform 1 0 1620 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1959
timestamp 1681620392
transform 1 0 1636 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1960
timestamp 1681620392
transform 1 0 1652 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1961
timestamp 1681620392
transform 1 0 1660 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2053
timestamp 1681620392
transform 1 0 1628 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1757
timestamp 1681620392
transform 1 0 1620 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1700
timestamp 1681620392
transform 1 0 1660 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1589
timestamp 1681620392
transform 1 0 1764 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1641
timestamp 1681620392
transform 1 0 1732 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1962
timestamp 1681620392
transform 1 0 1684 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1963
timestamp 1681620392
transform 1 0 1772 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1964
timestamp 1681620392
transform 1 0 1788 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1965
timestamp 1681620392
transform 1 0 1804 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1966
timestamp 1681620392
transform 1 0 1812 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2054
timestamp 1681620392
transform 1 0 1668 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2055
timestamp 1681620392
transform 1 0 1732 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1701
timestamp 1681620392
transform 1 0 1748 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2056
timestamp 1681620392
transform 1 0 1764 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1702
timestamp 1681620392
transform 1 0 1772 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2057
timestamp 1681620392
transform 1 0 1780 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2058
timestamp 1681620392
transform 1 0 1796 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2059
timestamp 1681620392
transform 1 0 1812 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1773
timestamp 1681620392
transform 1 0 1724 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1730
timestamp 1681620392
transform 1 0 1796 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1758
timestamp 1681620392
transform 1 0 1804 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1590
timestamp 1681620392
transform 1 0 1844 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1642
timestamp 1681620392
transform 1 0 1836 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1967
timestamp 1681620392
transform 1 0 1836 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1968
timestamp 1681620392
transform 1 0 1844 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1678
timestamp 1681620392
transform 1 0 1860 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_2060
timestamp 1681620392
transform 1 0 1860 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1643
timestamp 1681620392
transform 1 0 1884 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_2061
timestamp 1681620392
transform 1 0 1876 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2111
timestamp 1681620392
transform 1 0 1868 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_1613
timestamp 1681620392
transform 1 0 1948 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1644
timestamp 1681620392
transform 1 0 1916 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1969
timestamp 1681620392
transform 1 0 1908 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1970
timestamp 1681620392
transform 1 0 1916 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1679
timestamp 1681620392
transform 1 0 1924 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1971
timestamp 1681620392
transform 1 0 1932 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1972
timestamp 1681620392
transform 1 0 1948 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1703
timestamp 1681620392
transform 1 0 1916 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2062
timestamp 1681620392
transform 1 0 1924 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2063
timestamp 1681620392
transform 1 0 1940 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1731
timestamp 1681620392
transform 1 0 1924 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1732
timestamp 1681620392
transform 1 0 1940 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1645
timestamp 1681620392
transform 1 0 1996 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1973
timestamp 1681620392
transform 1 0 1980 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1680
timestamp 1681620392
transform 1 0 1988 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1974
timestamp 1681620392
transform 1 0 1996 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2064
timestamp 1681620392
transform 1 0 1988 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1704
timestamp 1681620392
transform 1 0 1996 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2065
timestamp 1681620392
transform 1 0 2004 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2066
timestamp 1681620392
transform 1 0 2020 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1733
timestamp 1681620392
transform 1 0 1988 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1734
timestamp 1681620392
transform 1 0 2004 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1787
timestamp 1681620392
transform 1 0 1980 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1759
timestamp 1681620392
transform 1 0 2020 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1646
timestamp 1681620392
transform 1 0 2068 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1647
timestamp 1681620392
transform 1 0 2092 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1648
timestamp 1681620392
transform 1 0 2132 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1649
timestamp 1681620392
transform 1 0 2164 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1650
timestamp 1681620392
transform 1 0 2204 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1975
timestamp 1681620392
transform 1 0 2116 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1976
timestamp 1681620392
transform 1 0 2132 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1977
timestamp 1681620392
transform 1 0 2148 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1978
timestamp 1681620392
transform 1 0 2164 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1979
timestamp 1681620392
transform 1 0 2172 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2067
timestamp 1681620392
transform 1 0 2068 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1705
timestamp 1681620392
transform 1 0 2132 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1681
timestamp 1681620392
transform 1 0 2180 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1651
timestamp 1681620392
transform 1 0 2244 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1980
timestamp 1681620392
transform 1 0 2188 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1981
timestamp 1681620392
transform 1 0 2204 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1982
timestamp 1681620392
transform 1 0 2212 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1983
timestamp 1681620392
transform 1 0 2228 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1984
timestamp 1681620392
transform 1 0 2244 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2068
timestamp 1681620392
transform 1 0 2140 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2069
timestamp 1681620392
transform 1 0 2164 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2070
timestamp 1681620392
transform 1 0 2180 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2071
timestamp 1681620392
transform 1 0 2196 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1735
timestamp 1681620392
transform 1 0 2164 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1736
timestamp 1681620392
transform 1 0 2188 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1760
timestamp 1681620392
transform 1 0 2172 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1774
timestamp 1681620392
transform 1 0 2156 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_2072
timestamp 1681620392
transform 1 0 2220 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2073
timestamp 1681620392
transform 1 0 2284 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1788
timestamp 1681620392
transform 1 0 2284 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1591
timestamp 1681620392
transform 1 0 2308 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1614
timestamp 1681620392
transform 1 0 2300 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1652
timestamp 1681620392
transform 1 0 2316 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1985
timestamp 1681620392
transform 1 0 2292 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1986
timestamp 1681620392
transform 1 0 2300 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1987
timestamp 1681620392
transform 1 0 2316 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1682
timestamp 1681620392
transform 1 0 2324 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1592
timestamp 1681620392
transform 1 0 2348 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1615
timestamp 1681620392
transform 1 0 2428 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1653
timestamp 1681620392
transform 1 0 2372 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1988
timestamp 1681620392
transform 1 0 2332 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1989
timestamp 1681620392
transform 1 0 2348 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2074
timestamp 1681620392
transform 1 0 2308 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2075
timestamp 1681620392
transform 1 0 2324 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1737
timestamp 1681620392
transform 1 0 2324 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1789
timestamp 1681620392
transform 1 0 2300 0 1 1885
box -3 -3 3 3
use M2_M1  M2_M1_2076
timestamp 1681620392
transform 1 0 2372 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1706
timestamp 1681620392
transform 1 0 2412 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1654
timestamp 1681620392
transform 1 0 2444 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1990
timestamp 1681620392
transform 1 0 2452 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2077
timestamp 1681620392
transform 1 0 2444 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1707
timestamp 1681620392
transform 1 0 2452 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1738
timestamp 1681620392
transform 1 0 2444 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1655
timestamp 1681620392
transform 1 0 2476 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1991
timestamp 1681620392
transform 1 0 2476 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2078
timestamp 1681620392
transform 1 0 2476 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1992
timestamp 1681620392
transform 1 0 2500 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1708
timestamp 1681620392
transform 1 0 2500 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2079
timestamp 1681620392
transform 1 0 2508 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2112
timestamp 1681620392
transform 1 0 2508 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_1616
timestamp 1681620392
transform 1 0 2540 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1656
timestamp 1681620392
transform 1 0 2540 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1683
timestamp 1681620392
transform 1 0 2532 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1993
timestamp 1681620392
transform 1 0 2540 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2080
timestamp 1681620392
transform 1 0 2532 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1790
timestamp 1681620392
transform 1 0 2524 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1739
timestamp 1681620392
transform 1 0 2540 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1657
timestamp 1681620392
transform 1 0 2636 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1994
timestamp 1681620392
transform 1 0 2556 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2081
timestamp 1681620392
transform 1 0 2580 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2082
timestamp 1681620392
transform 1 0 2636 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1740
timestamp 1681620392
transform 1 0 2580 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1791
timestamp 1681620392
transform 1 0 2564 0 1 1885
box -3 -3 3 3
use M2_M1  M2_M1_1995
timestamp 1681620392
transform 1 0 2668 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1617
timestamp 1681620392
transform 1 0 2716 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1658
timestamp 1681620392
transform 1 0 2708 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1684
timestamp 1681620392
transform 1 0 2684 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1685
timestamp 1681620392
transform 1 0 2700 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_1996
timestamp 1681620392
transform 1 0 2708 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1997
timestamp 1681620392
transform 1 0 2716 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1709
timestamp 1681620392
transform 1 0 2676 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2113
timestamp 1681620392
transform 1 0 2676 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2083
timestamp 1681620392
transform 1 0 2700 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1593
timestamp 1681620392
transform 1 0 2740 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1618
timestamp 1681620392
transform 1 0 2740 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1659
timestamp 1681620392
transform 1 0 2732 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_1998
timestamp 1681620392
transform 1 0 2732 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2084
timestamp 1681620392
transform 1 0 2724 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1741
timestamp 1681620392
transform 1 0 2716 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1761
timestamp 1681620392
transform 1 0 2716 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1762
timestamp 1681620392
transform 1 0 2740 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1710
timestamp 1681620392
transform 1 0 2748 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1594
timestamp 1681620392
transform 1 0 2836 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1619
timestamp 1681620392
transform 1 0 2788 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1620
timestamp 1681620392
transform 1 0 2828 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1660
timestamp 1681620392
transform 1 0 2828 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1595
timestamp 1681620392
transform 1 0 2900 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_1999
timestamp 1681620392
transform 1 0 2788 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2000
timestamp 1681620392
transform 1 0 2876 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2001
timestamp 1681620392
transform 1 0 2892 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2085
timestamp 1681620392
transform 1 0 2772 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2086
timestamp 1681620392
transform 1 0 2780 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2087
timestamp 1681620392
transform 1 0 2788 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2088
timestamp 1681620392
transform 1 0 2852 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2114
timestamp 1681620392
transform 1 0 2772 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_1742
timestamp 1681620392
transform 1 0 2780 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1743
timestamp 1681620392
transform 1 0 2796 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1763
timestamp 1681620392
transform 1 0 2876 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1661
timestamp 1681620392
transform 1 0 2916 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1662
timestamp 1681620392
transform 1 0 2956 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_2002
timestamp 1681620392
transform 1 0 2916 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2003
timestamp 1681620392
transform 1 0 2932 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_1686
timestamp 1681620392
transform 1 0 3012 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_2089
timestamp 1681620392
transform 1 0 2900 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1711
timestamp 1681620392
transform 1 0 2916 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2090
timestamp 1681620392
transform 1 0 2956 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_1712
timestamp 1681620392
transform 1 0 2996 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_2091
timestamp 1681620392
transform 1 0 3012 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2115
timestamp 1681620392
transform 1 0 2916 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_1744
timestamp 1681620392
transform 1 0 3028 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1764
timestamp 1681620392
transform 1 0 2932 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1792
timestamp 1681620392
transform 1 0 3028 0 1 1885
box -3 -3 3 3
use Project_Top_VIA0  Project_Top_VIA0_22
timestamp 1681620392
transform 1 0 24 0 1 1870
box -10 -3 10 3
use FILL  FILL_367
timestamp 1681620392
transform 1 0 72 0 -1 1970
box -8 -3 16 105
use FILL  FILL_368
timestamp 1681620392
transform 1 0 80 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_23
timestamp 1681620392
transform 1 0 88 0 -1 1970
box -8 -3 46 105
use FILL  FILL_369
timestamp 1681620392
transform 1 0 128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_370
timestamp 1681620392
transform 1 0 136 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_24
timestamp 1681620392
transform 1 0 144 0 -1 1970
box -8 -3 46 105
use FILL  FILL_371
timestamp 1681620392
transform 1 0 184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_372
timestamp 1681620392
transform 1 0 192 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_105
timestamp 1681620392
transform -1 0 216 0 -1 1970
box -9 -3 26 105
use NOR2X1  NOR2X1_31
timestamp 1681620392
transform 1 0 216 0 -1 1970
box -8 -3 32 105
use FILL  FILL_374
timestamp 1681620392
transform 1 0 240 0 -1 1970
box -8 -3 16 105
use FILL  FILL_376
timestamp 1681620392
transform 1 0 248 0 -1 1970
box -8 -3 16 105
use FILL  FILL_378
timestamp 1681620392
transform 1 0 256 0 -1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_35
timestamp 1681620392
transform 1 0 264 0 -1 1970
box -8 -3 32 105
use OAI22X1  OAI22X1_8
timestamp 1681620392
transform 1 0 288 0 -1 1970
box -8 -3 46 105
use AOI21X1  AOI21X1_9
timestamp 1681620392
transform -1 0 360 0 -1 1970
box -7 -3 39 105
use INVX2  INVX2_116
timestamp 1681620392
transform 1 0 360 0 -1 1970
box -9 -3 26 105
use NAND3X1  NAND3X1_41
timestamp 1681620392
transform 1 0 376 0 -1 1970
box -8 -3 40 105
use OAI21X1  OAI21X1_127
timestamp 1681620392
transform -1 0 440 0 -1 1970
box -8 -3 34 105
use OR2X2  OR2X2_1
timestamp 1681620392
transform 1 0 440 0 -1 1970
box -7 -3 35 105
use NAND2X1  NAND2X1_112
timestamp 1681620392
transform -1 0 496 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_113
timestamp 1681620392
transform -1 0 520 0 -1 1970
box -8 -3 32 105
use OAI22X1  OAI22X1_9
timestamp 1681620392
transform -1 0 560 0 -1 1970
box -8 -3 46 105
use NOR2X1  NOR2X1_36
timestamp 1681620392
transform 1 0 560 0 -1 1970
box -8 -3 32 105
use INVX2  INVX2_117
timestamp 1681620392
transform 1 0 584 0 -1 1970
box -9 -3 26 105
use OAI21X1  OAI21X1_128
timestamp 1681620392
transform 1 0 600 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_129
timestamp 1681620392
transform -1 0 664 0 -1 1970
box -8 -3 34 105
use M3_M2  M3_M2_1793
timestamp 1681620392
transform 1 0 692 0 1 1875
box -3 -3 3 3
use INVX2  INVX2_118
timestamp 1681620392
transform 1 0 664 0 -1 1970
box -9 -3 26 105
use OR2X1  OR2X1_5
timestamp 1681620392
transform 1 0 680 0 -1 1970
box -8 -3 40 105
use BUFX2  BUFX2_14
timestamp 1681620392
transform -1 0 736 0 -1 1970
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_121
timestamp 1681620392
transform -1 0 832 0 -1 1970
box -8 -3 104 105
use NOR2X1  NOR2X1_37
timestamp 1681620392
transform 1 0 832 0 -1 1970
box -8 -3 32 105
use INVX2  INVX2_119
timestamp 1681620392
transform 1 0 856 0 -1 1970
box -9 -3 26 105
use NAND3X1  NAND3X1_42
timestamp 1681620392
transform 1 0 872 0 -1 1970
box -8 -3 40 105
use FILL  FILL_404
timestamp 1681620392
transform 1 0 904 0 -1 1970
box -8 -3 16 105
use FILL  FILL_405
timestamp 1681620392
transform 1 0 912 0 -1 1970
box -8 -3 16 105
use FILL  FILL_406
timestamp 1681620392
transform 1 0 920 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_10
timestamp 1681620392
transform -1 0 968 0 -1 1970
box -8 -3 46 105
use FILL  FILL_407
timestamp 1681620392
transform 1 0 968 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_11
timestamp 1681620392
transform -1 0 1016 0 -1 1970
box -8 -3 46 105
use FILL  FILL_408
timestamp 1681620392
transform 1 0 1016 0 -1 1970
box -8 -3 16 105
use FILL  FILL_409
timestamp 1681620392
transform 1 0 1024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_410
timestamp 1681620392
transform 1 0 1032 0 -1 1970
box -8 -3 16 105
use FILL  FILL_411
timestamp 1681620392
transform 1 0 1040 0 -1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_43
timestamp 1681620392
transform -1 0 1080 0 -1 1970
box -8 -3 40 105
use FILL  FILL_412
timestamp 1681620392
transform 1 0 1080 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_120
timestamp 1681620392
transform 1 0 1088 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_121
timestamp 1681620392
transform 1 0 1104 0 -1 1970
box -9 -3 26 105
use FILL  FILL_413
timestamp 1681620392
transform 1 0 1120 0 -1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_44
timestamp 1681620392
transform 1 0 1128 0 -1 1970
box -8 -3 40 105
use INVX2  INVX2_122
timestamp 1681620392
transform 1 0 1160 0 -1 1970
box -9 -3 26 105
use M3_M2  M3_M2_1794
timestamp 1681620392
transform 1 0 1212 0 1 1875
box -3 -3 3 3
use NAND3X1  NAND3X1_45
timestamp 1681620392
transform 1 0 1176 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_46
timestamp 1681620392
transform 1 0 1208 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_47
timestamp 1681620392
transform -1 0 1272 0 -1 1970
box -8 -3 40 105
use M3_M2  M3_M2_1795
timestamp 1681620392
transform 1 0 1372 0 1 1875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_122
timestamp 1681620392
transform -1 0 1368 0 -1 1970
box -8 -3 104 105
use FILL  FILL_414
timestamp 1681620392
transform 1 0 1368 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_1796
timestamp 1681620392
transform 1 0 1444 0 1 1875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_123
timestamp 1681620392
transform 1 0 1376 0 -1 1970
box -8 -3 104 105
use FILL  FILL_415
timestamp 1681620392
transform 1 0 1472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_416
timestamp 1681620392
transform 1 0 1480 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_123
timestamp 1681620392
transform 1 0 1488 0 -1 1970
box -9 -3 26 105
use FILL  FILL_417
timestamp 1681620392
transform 1 0 1504 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_124
timestamp 1681620392
transform -1 0 1528 0 -1 1970
box -9 -3 26 105
use FILL  FILL_418
timestamp 1681620392
transform 1 0 1528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_419
timestamp 1681620392
transform 1 0 1536 0 -1 1970
box -8 -3 16 105
use FILL  FILL_420
timestamp 1681620392
transform 1 0 1544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_422
timestamp 1681620392
transform 1 0 1552 0 -1 1970
box -8 -3 16 105
use FILL  FILL_423
timestamp 1681620392
transform 1 0 1560 0 -1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_131
timestamp 1681620392
transform -1 0 1600 0 -1 1970
box -8 -3 34 105
use FILL  FILL_424
timestamp 1681620392
transform 1 0 1600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_434
timestamp 1681620392
transform 1 0 1608 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_14
timestamp 1681620392
transform -1 0 1656 0 -1 1970
box -8 -3 46 105
use INVX2  INVX2_129
timestamp 1681620392
transform 1 0 1656 0 -1 1970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_130
timestamp 1681620392
transform 1 0 1672 0 -1 1970
box -8 -3 104 105
use OAI22X1  OAI22X1_15
timestamp 1681620392
transform 1 0 1768 0 -1 1970
box -8 -3 46 105
use OAI21X1  OAI21X1_136
timestamp 1681620392
transform 1 0 1808 0 -1 1970
box -8 -3 34 105
use NAND2X1  NAND2X1_115
timestamp 1681620392
transform 1 0 1840 0 -1 1970
box -8 -3 32 105
use FILL  FILL_435
timestamp 1681620392
transform 1 0 1864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_436
timestamp 1681620392
transform 1 0 1872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_437
timestamp 1681620392
transform 1 0 1880 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_15
timestamp 1681620392
transform 1 0 1888 0 -1 1970
box -5 -3 28 105
use OAI22X1  OAI22X1_16
timestamp 1681620392
transform 1 0 1912 0 -1 1970
box -8 -3 46 105
use FILL  FILL_438
timestamp 1681620392
transform 1 0 1952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_439
timestamp 1681620392
transform 1 0 1960 0 -1 1970
box -8 -3 16 105
use FILL  FILL_440
timestamp 1681620392
transform 1 0 1968 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_17
timestamp 1681620392
transform -1 0 2016 0 -1 1970
box -8 -3 46 105
use INVX2  INVX2_130
timestamp 1681620392
transform -1 0 2032 0 -1 1970
box -9 -3 26 105
use M3_M2  M3_M2_1797
timestamp 1681620392
transform 1 0 2092 0 1 1875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_131
timestamp 1681620392
transform -1 0 2128 0 -1 1970
box -8 -3 104 105
use OAI22X1  OAI22X1_18
timestamp 1681620392
transform -1 0 2168 0 -1 1970
box -8 -3 46 105
use M3_M2  M3_M2_1798
timestamp 1681620392
transform 1 0 2196 0 1 1875
box -3 -3 3 3
use OAI22X1  OAI22X1_19
timestamp 1681620392
transform -1 0 2208 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_20
timestamp 1681620392
transform -1 0 2248 0 -1 1970
box -8 -3 46 105
use INVX2  INVX2_131
timestamp 1681620392
transform -1 0 2264 0 -1 1970
box -9 -3 26 105
use FILL  FILL_441
timestamp 1681620392
transform 1 0 2264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_442
timestamp 1681620392
transform 1 0 2272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_443
timestamp 1681620392
transform 1 0 2280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_444
timestamp 1681620392
transform 1 0 2288 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_21
timestamp 1681620392
transform -1 0 2336 0 -1 1970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_132
timestamp 1681620392
transform 1 0 2336 0 -1 1970
box -8 -3 104 105
use INVX2  INVX2_132
timestamp 1681620392
transform 1 0 2432 0 -1 1970
box -9 -3 26 105
use FILL  FILL_445
timestamp 1681620392
transform 1 0 2448 0 -1 1970
box -8 -3 16 105
use FILL  FILL_446
timestamp 1681620392
transform 1 0 2456 0 -1 1970
box -8 -3 16 105
use FILL  FILL_447
timestamp 1681620392
transform 1 0 2464 0 -1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_137
timestamp 1681620392
transform 1 0 2472 0 -1 1970
box -8 -3 34 105
use NAND2X1  NAND2X1_116
timestamp 1681620392
transform -1 0 2528 0 -1 1970
box -8 -3 32 105
use FILL  FILL_448
timestamp 1681620392
transform 1 0 2528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_450
timestamp 1681620392
transform 1 0 2536 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_134
timestamp 1681620392
transform 1 0 2544 0 -1 1970
box -8 -3 104 105
use FILL  FILL_453
timestamp 1681620392
transform 1 0 2640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_454
timestamp 1681620392
transform 1 0 2648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_456
timestamp 1681620392
transform 1 0 2656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_458
timestamp 1681620392
transform 1 0 2664 0 -1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_142
timestamp 1681620392
transform -1 0 2704 0 -1 1970
box -8 -3 34 105
use FILL  FILL_459
timestamp 1681620392
transform 1 0 2704 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_136
timestamp 1681620392
transform 1 0 2712 0 -1 1970
box -9 -3 26 105
use FILL  FILL_460
timestamp 1681620392
transform 1 0 2728 0 -1 1970
box -8 -3 16 105
use FILL  FILL_461
timestamp 1681620392
transform 1 0 2736 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_1799
timestamp 1681620392
transform 1 0 2756 0 1 1875
box -3 -3 3 3
use FILL  FILL_462
timestamp 1681620392
transform 1 0 2744 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_137
timestamp 1681620392
transform 1 0 2752 0 -1 1970
box -9 -3 26 105
use M3_M2  M3_M2_1800
timestamp 1681620392
transform 1 0 2788 0 1 1875
box -3 -3 3 3
use NAND2X1  NAND2X1_119
timestamp 1681620392
transform -1 0 2792 0 -1 1970
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_136
timestamp 1681620392
transform -1 0 2888 0 -1 1970
box -8 -3 104 105
use OAI21X1  OAI21X1_143
timestamp 1681620392
transform 1 0 2888 0 -1 1970
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_137
timestamp 1681620392
transform 1 0 2920 0 -1 1970
box -8 -3 104 105
use Project_Top_VIA0  Project_Top_VIA0_23
timestamp 1681620392
transform 1 0 3067 0 1 1870
box -10 -3 10 3
use M3_M2  M3_M2_1855
timestamp 1681620392
transform 1 0 92 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_2127
timestamp 1681620392
transform 1 0 108 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2161
timestamp 1681620392
transform 1 0 92 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2162
timestamp 1681620392
transform 1 0 108 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2257
timestamp 1681620392
transform 1 0 84 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1908
timestamp 1681620392
transform 1 0 100 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_2258
timestamp 1681620392
transform 1 0 108 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1856
timestamp 1681620392
transform 1 0 124 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_2163
timestamp 1681620392
transform 1 0 124 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2259
timestamp 1681620392
transform 1 0 140 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2260
timestamp 1681620392
transform 1 0 148 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1924
timestamp 1681620392
transform 1 0 140 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_2128
timestamp 1681620392
transform 1 0 172 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2164
timestamp 1681620392
transform 1 0 204 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2261
timestamp 1681620392
transform 1 0 172 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1909
timestamp 1681620392
transform 1 0 180 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_2262
timestamp 1681620392
transform 1 0 188 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1925
timestamp 1681620392
transform 1 0 164 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1952
timestamp 1681620392
transform 1 0 148 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_2344
timestamp 1681620392
transform 1 0 180 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_2165
timestamp 1681620392
transform 1 0 228 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2263
timestamp 1681620392
transform 1 0 212 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2345
timestamp 1681620392
transform 1 0 220 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_1953
timestamp 1681620392
transform 1 0 220 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_2166
timestamp 1681620392
transform 1 0 244 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1954
timestamp 1681620392
transform 1 0 244 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1811
timestamp 1681620392
transform 1 0 324 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1826
timestamp 1681620392
transform 1 0 308 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1827
timestamp 1681620392
transform 1 0 324 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_2129
timestamp 1681620392
transform 1 0 292 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2130
timestamp 1681620392
transform 1 0 316 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2131
timestamp 1681620392
transform 1 0 324 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2167
timestamp 1681620392
transform 1 0 284 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2264
timestamp 1681620392
transform 1 0 268 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2265
timestamp 1681620392
transform 1 0 276 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2168
timestamp 1681620392
transform 1 0 324 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2266
timestamp 1681620392
transform 1 0 300 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2267
timestamp 1681620392
transform 1 0 316 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1926
timestamp 1681620392
transform 1 0 300 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1818
timestamp 1681620392
transform 1 0 348 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1882
timestamp 1681620392
transform 1 0 356 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_2268
timestamp 1681620392
transform 1 0 348 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2269
timestamp 1681620392
transform 1 0 356 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1927
timestamp 1681620392
transform 1 0 356 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_2132
timestamp 1681620392
transform 1 0 380 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1883
timestamp 1681620392
transform 1 0 380 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1828
timestamp 1681620392
transform 1 0 396 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1829
timestamp 1681620392
transform 1 0 420 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_2133
timestamp 1681620392
transform 1 0 396 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2169
timestamp 1681620392
transform 1 0 388 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2270
timestamp 1681620392
transform 1 0 380 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1857
timestamp 1681620392
transform 1 0 412 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_2134
timestamp 1681620392
transform 1 0 420 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2135
timestamp 1681620392
transform 1 0 428 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2170
timestamp 1681620392
transform 1 0 412 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2271
timestamp 1681620392
transform 1 0 404 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1884
timestamp 1681620392
transform 1 0 428 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1812
timestamp 1681620392
transform 1 0 476 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1819
timestamp 1681620392
transform 1 0 484 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1858
timestamp 1681620392
transform 1 0 444 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1859
timestamp 1681620392
transform 1 0 468 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_2136
timestamp 1681620392
transform 1 0 476 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2171
timestamp 1681620392
transform 1 0 436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2172
timestamp 1681620392
transform 1 0 444 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1910
timestamp 1681620392
transform 1 0 420 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_2272
timestamp 1681620392
transform 1 0 444 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2273
timestamp 1681620392
transform 1 0 452 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1928
timestamp 1681620392
transform 1 0 444 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_2173
timestamp 1681620392
transform 1 0 476 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1830
timestamp 1681620392
transform 1 0 508 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_2137
timestamp 1681620392
transform 1 0 500 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1885
timestamp 1681620392
transform 1 0 500 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_2274
timestamp 1681620392
transform 1 0 476 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2275
timestamp 1681620392
transform 1 0 484 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2276
timestamp 1681620392
transform 1 0 500 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1929
timestamp 1681620392
transform 1 0 492 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_2346
timestamp 1681620392
transform 1 0 508 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_1955
timestamp 1681620392
transform 1 0 484 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1956
timestamp 1681620392
transform 1 0 500 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1831
timestamp 1681620392
transform 1 0 532 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1813
timestamp 1681620392
transform 1 0 628 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_2174
timestamp 1681620392
transform 1 0 524 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2175
timestamp 1681620392
transform 1 0 580 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1886
timestamp 1681620392
transform 1 0 588 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_2176
timestamp 1681620392
transform 1 0 620 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2177
timestamp 1681620392
transform 1 0 636 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2178
timestamp 1681620392
transform 1 0 652 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2277
timestamp 1681620392
transform 1 0 540 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1911
timestamp 1681620392
transform 1 0 588 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_2278
timestamp 1681620392
transform 1 0 628 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2279
timestamp 1681620392
transform 1 0 644 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1957
timestamp 1681620392
transform 1 0 540 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1912
timestamp 1681620392
transform 1 0 652 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1860
timestamp 1681620392
transform 1 0 740 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1814
timestamp 1681620392
transform 1 0 868 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1832
timestamp 1681620392
transform 1 0 820 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1861
timestamp 1681620392
transform 1 0 868 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_2138
timestamp 1681620392
transform 1 0 876 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2179
timestamp 1681620392
transform 1 0 700 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2180
timestamp 1681620392
transform 1 0 764 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2181
timestamp 1681620392
transform 1 0 772 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1887
timestamp 1681620392
transform 1 0 788 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_2182
timestamp 1681620392
transform 1 0 836 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2183
timestamp 1681620392
transform 1 0 876 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2280
timestamp 1681620392
transform 1 0 660 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2281
timestamp 1681620392
transform 1 0 676 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2282
timestamp 1681620392
transform 1 0 764 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1930
timestamp 1681620392
transform 1 0 644 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1931
timestamp 1681620392
transform 1 0 700 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1958
timestamp 1681620392
transform 1 0 676 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1959
timestamp 1681620392
transform 1 0 700 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_2283
timestamp 1681620392
transform 1 0 788 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1932
timestamp 1681620392
transform 1 0 836 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1960
timestamp 1681620392
transform 1 0 772 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1833
timestamp 1681620392
transform 1 0 892 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_2123
timestamp 1681620392
transform 1 0 924 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_2139
timestamp 1681620392
transform 1 0 892 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2140
timestamp 1681620392
transform 1 0 916 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2141
timestamp 1681620392
transform 1 0 932 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2184
timestamp 1681620392
transform 1 0 892 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2185
timestamp 1681620392
transform 1 0 916 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2284
timestamp 1681620392
transform 1 0 892 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2186
timestamp 1681620392
transform 1 0 940 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2187
timestamp 1681620392
transform 1 0 956 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2188
timestamp 1681620392
transform 1 0 964 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2285
timestamp 1681620392
transform 1 0 932 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1961
timestamp 1681620392
transform 1 0 916 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1962
timestamp 1681620392
transform 1 0 932 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1913
timestamp 1681620392
transform 1 0 964 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1815
timestamp 1681620392
transform 1 0 988 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1801
timestamp 1681620392
transform 1 0 1148 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1820
timestamp 1681620392
transform 1 0 1124 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1834
timestamp 1681620392
transform 1 0 1012 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1835
timestamp 1681620392
transform 1 0 1076 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1836
timestamp 1681620392
transform 1 0 1116 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1821
timestamp 1681620392
transform 1 0 1164 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_2124
timestamp 1681620392
transform 1 0 1124 0 1 1835
box -2 -2 2 2
use M3_M2  M3_M2_1862
timestamp 1681620392
transform 1 0 996 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1863
timestamp 1681620392
transform 1 0 1052 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_2142
timestamp 1681620392
transform 1 0 1116 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2189
timestamp 1681620392
transform 1 0 988 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2190
timestamp 1681620392
transform 1 0 1012 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2191
timestamp 1681620392
transform 1 0 1020 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2192
timestamp 1681620392
transform 1 0 1052 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2286
timestamp 1681620392
transform 1 0 980 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2287
timestamp 1681620392
transform 1 0 996 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1914
timestamp 1681620392
transform 1 0 1004 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1888
timestamp 1681620392
transform 1 0 1100 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_2288
timestamp 1681620392
transform 1 0 1012 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2289
timestamp 1681620392
transform 1 0 1100 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1933
timestamp 1681620392
transform 1 0 996 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1934
timestamp 1681620392
transform 1 0 1100 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1837
timestamp 1681620392
transform 1 0 1148 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_2125
timestamp 1681620392
transform 1 0 1180 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_2143
timestamp 1681620392
transform 1 0 1140 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2144
timestamp 1681620392
transform 1 0 1164 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2193
timestamp 1681620392
transform 1 0 1124 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1889
timestamp 1681620392
transform 1 0 1132 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_2194
timestamp 1681620392
transform 1 0 1148 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1915
timestamp 1681620392
transform 1 0 1132 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1890
timestamp 1681620392
transform 1 0 1164 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1802
timestamp 1681620392
transform 1 0 1212 0 1 1865
box -3 -3 3 3
use M2_M1  M2_M1_2145
timestamp 1681620392
transform 1 0 1188 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2195
timestamp 1681620392
transform 1 0 1172 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2290
timestamp 1681620392
transform 1 0 1148 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1891
timestamp 1681620392
transform 1 0 1204 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_2196
timestamp 1681620392
transform 1 0 1228 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1892
timestamp 1681620392
transform 1 0 1252 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1893
timestamp 1681620392
transform 1 0 1268 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1864
timestamp 1681620392
transform 1 0 1300 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_2146
timestamp 1681620392
transform 1 0 1308 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1865
timestamp 1681620392
transform 1 0 1332 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1803
timestamp 1681620392
transform 1 0 1372 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1838
timestamp 1681620392
transform 1 0 1364 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_2197
timestamp 1681620392
transform 1 0 1284 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2198
timestamp 1681620392
transform 1 0 1300 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2199
timestamp 1681620392
transform 1 0 1308 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2200
timestamp 1681620392
transform 1 0 1332 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2201
timestamp 1681620392
transform 1 0 1348 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2291
timestamp 1681620392
transform 1 0 1204 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1916
timestamp 1681620392
transform 1 0 1228 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_2292
timestamp 1681620392
transform 1 0 1292 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1935
timestamp 1681620392
transform 1 0 1204 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1963
timestamp 1681620392
transform 1 0 1228 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1894
timestamp 1681620392
transform 1 0 1356 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_2202
timestamp 1681620392
transform 1 0 1372 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2293
timestamp 1681620392
transform 1 0 1348 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2294
timestamp 1681620392
transform 1 0 1356 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2295
timestamp 1681620392
transform 1 0 1364 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1964
timestamp 1681620392
transform 1 0 1340 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_2347
timestamp 1681620392
transform 1 0 1364 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_2203
timestamp 1681620392
transform 1 0 1396 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1839
timestamp 1681620392
transform 1 0 1428 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1866
timestamp 1681620392
transform 1 0 1436 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1867
timestamp 1681620392
transform 1 0 1460 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1804
timestamp 1681620392
transform 1 0 1532 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1840
timestamp 1681620392
transform 1 0 1500 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_2147
timestamp 1681620392
transform 1 0 1484 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2204
timestamp 1681620392
transform 1 0 1428 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2205
timestamp 1681620392
transform 1 0 1436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2296
timestamp 1681620392
transform 1 0 1420 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1895
timestamp 1681620392
transform 1 0 1452 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_2206
timestamp 1681620392
transform 1 0 1468 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1896
timestamp 1681620392
transform 1 0 1484 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1868
timestamp 1681620392
transform 1 0 1524 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1841
timestamp 1681620392
transform 1 0 1556 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1869
timestamp 1681620392
transform 1 0 1572 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_2207
timestamp 1681620392
transform 1 0 1500 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2208
timestamp 1681620392
transform 1 0 1516 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2209
timestamp 1681620392
transform 1 0 1524 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2210
timestamp 1681620392
transform 1 0 1540 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2211
timestamp 1681620392
transform 1 0 1556 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2297
timestamp 1681620392
transform 1 0 1452 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2298
timestamp 1681620392
transform 1 0 1460 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2299
timestamp 1681620392
transform 1 0 1484 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2300
timestamp 1681620392
transform 1 0 1492 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2301
timestamp 1681620392
transform 1 0 1508 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2302
timestamp 1681620392
transform 1 0 1524 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2303
timestamp 1681620392
transform 1 0 1548 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1936
timestamp 1681620392
transform 1 0 1516 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1937
timestamp 1681620392
transform 1 0 1532 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1897
timestamp 1681620392
transform 1 0 1564 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_2148
timestamp 1681620392
transform 1 0 1588 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1822
timestamp 1681620392
transform 1 0 1692 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_2212
timestamp 1681620392
transform 1 0 1580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2213
timestamp 1681620392
transform 1 0 1596 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2304
timestamp 1681620392
transform 1 0 1564 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2305
timestamp 1681620392
transform 1 0 1572 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1938
timestamp 1681620392
transform 1 0 1564 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1898
timestamp 1681620392
transform 1 0 1604 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_2214
timestamp 1681620392
transform 1 0 1636 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1805
timestamp 1681620392
transform 1 0 1716 0 1 1865
box -3 -3 3 3
use M2_M1  M2_M1_2149
timestamp 1681620392
transform 1 0 1716 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2215
timestamp 1681620392
transform 1 0 1700 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2306
timestamp 1681620392
transform 1 0 1676 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2307
timestamp 1681620392
transform 1 0 1692 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2308
timestamp 1681620392
transform 1 0 1716 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2309
timestamp 1681620392
transform 1 0 1724 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1939
timestamp 1681620392
transform 1 0 1724 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1965
timestamp 1681620392
transform 1 0 1716 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1842
timestamp 1681620392
transform 1 0 1764 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1870
timestamp 1681620392
transform 1 0 1748 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1899
timestamp 1681620392
transform 1 0 1740 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1823
timestamp 1681620392
transform 1 0 1788 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1843
timestamp 1681620392
transform 1 0 1860 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1871
timestamp 1681620392
transform 1 0 1812 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_2216
timestamp 1681620392
transform 1 0 1748 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2217
timestamp 1681620392
transform 1 0 1764 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1900
timestamp 1681620392
transform 1 0 1772 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_2218
timestamp 1681620392
transform 1 0 1812 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2310
timestamp 1681620392
transform 1 0 1756 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2311
timestamp 1681620392
transform 1 0 1772 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2312
timestamp 1681620392
transform 1 0 1788 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1940
timestamp 1681620392
transform 1 0 1756 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1941
timestamp 1681620392
transform 1 0 1812 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1942
timestamp 1681620392
transform 1 0 1828 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1844
timestamp 1681620392
transform 1 0 1884 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1872
timestamp 1681620392
transform 1 0 1884 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_2219
timestamp 1681620392
transform 1 0 1884 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2150
timestamp 1681620392
transform 1 0 1908 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1901
timestamp 1681620392
transform 1 0 1908 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_2220
timestamp 1681620392
transform 1 0 1916 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2313
timestamp 1681620392
transform 1 0 1892 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1917
timestamp 1681620392
transform 1 0 1900 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_2314
timestamp 1681620392
transform 1 0 1908 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1943
timestamp 1681620392
transform 1 0 1892 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_2221
timestamp 1681620392
transform 1 0 1932 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1902
timestamp 1681620392
transform 1 0 1948 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_2222
timestamp 1681620392
transform 1 0 1956 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2315
timestamp 1681620392
transform 1 0 1940 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2316
timestamp 1681620392
transform 1 0 1956 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1944
timestamp 1681620392
transform 1 0 1956 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1873
timestamp 1681620392
transform 1 0 2028 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_2223
timestamp 1681620392
transform 1 0 2004 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1903
timestamp 1681620392
transform 1 0 2012 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_2224
timestamp 1681620392
transform 1 0 2028 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2317
timestamp 1681620392
transform 1 0 1988 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2318
timestamp 1681620392
transform 1 0 1996 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2319
timestamp 1681620392
transform 1 0 2012 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2320
timestamp 1681620392
transform 1 0 2028 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1945
timestamp 1681620392
transform 1 0 2028 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1806
timestamp 1681620392
transform 1 0 2052 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1845
timestamp 1681620392
transform 1 0 2060 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_2151
timestamp 1681620392
transform 1 0 2060 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1874
timestamp 1681620392
transform 1 0 2068 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_2225
timestamp 1681620392
transform 1 0 2052 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2226
timestamp 1681620392
transform 1 0 2068 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2321
timestamp 1681620392
transform 1 0 2044 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1918
timestamp 1681620392
transform 1 0 2052 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1919
timestamp 1681620392
transform 1 0 2068 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1807
timestamp 1681620392
transform 1 0 2140 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1808
timestamp 1681620392
transform 1 0 2180 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1875
timestamp 1681620392
transform 1 0 2124 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1904
timestamp 1681620392
transform 1 0 2092 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1905
timestamp 1681620392
transform 1 0 2116 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_2227
timestamp 1681620392
transform 1 0 2140 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2322
timestamp 1681620392
transform 1 0 2076 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2323
timestamp 1681620392
transform 1 0 2092 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1966
timestamp 1681620392
transform 1 0 2060 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1809
timestamp 1681620392
transform 1 0 2220 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1846
timestamp 1681620392
transform 1 0 2204 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_2228
timestamp 1681620392
transform 1 0 2188 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1876
timestamp 1681620392
transform 1 0 2212 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1810
timestamp 1681620392
transform 1 0 2308 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1847
timestamp 1681620392
transform 1 0 2340 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1877
timestamp 1681620392
transform 1 0 2324 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1848
timestamp 1681620392
transform 1 0 2372 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1878
timestamp 1681620392
transform 1 0 2468 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_2229
timestamp 1681620392
transform 1 0 2236 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2230
timestamp 1681620392
transform 1 0 2292 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2231
timestamp 1681620392
transform 1 0 2308 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2232
timestamp 1681620392
transform 1 0 2324 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2233
timestamp 1681620392
transform 1 0 2332 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2234
timestamp 1681620392
transform 1 0 2348 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2235
timestamp 1681620392
transform 1 0 2372 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2236
timestamp 1681620392
transform 1 0 2412 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2324
timestamp 1681620392
transform 1 0 2212 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2325
timestamp 1681620392
transform 1 0 2300 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1967
timestamp 1681620392
transform 1 0 2212 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1920
timestamp 1681620392
transform 1 0 2308 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_2326
timestamp 1681620392
transform 1 0 2316 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1921
timestamp 1681620392
transform 1 0 2332 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_2327
timestamp 1681620392
transform 1 0 2340 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1922
timestamp 1681620392
transform 1 0 2348 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_2328
timestamp 1681620392
transform 1 0 2356 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2329
timestamp 1681620392
transform 1 0 2372 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2330
timestamp 1681620392
transform 1 0 2388 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1946
timestamp 1681620392
transform 1 0 2316 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1947
timestamp 1681620392
transform 1 0 2412 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1968
timestamp 1681620392
transform 1 0 2388 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1849
timestamp 1681620392
transform 1 0 2492 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1879
timestamp 1681620392
transform 1 0 2484 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_2237
timestamp 1681620392
transform 1 0 2484 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2238
timestamp 1681620392
transform 1 0 2492 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2331
timestamp 1681620392
transform 1 0 2492 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1850
timestamp 1681620392
transform 1 0 2516 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_2152
timestamp 1681620392
transform 1 0 2532 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2239
timestamp 1681620392
transform 1 0 2508 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2240
timestamp 1681620392
transform 1 0 2516 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1923
timestamp 1681620392
transform 1 0 2516 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_2332
timestamp 1681620392
transform 1 0 2540 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2333
timestamp 1681620392
transform 1 0 2548 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2241
timestamp 1681620392
transform 1 0 2564 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2242
timestamp 1681620392
transform 1 0 2580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2153
timestamp 1681620392
transform 1 0 2604 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2334
timestamp 1681620392
transform 1 0 2604 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1851
timestamp 1681620392
transform 1 0 2620 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_2243
timestamp 1681620392
transform 1 0 2620 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1816
timestamp 1681620392
transform 1 0 2684 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_2244
timestamp 1681620392
transform 1 0 2668 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2335
timestamp 1681620392
transform 1 0 2652 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2336
timestamp 1681620392
transform 1 0 2660 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2348
timestamp 1681620392
transform 1 0 2636 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_1948
timestamp 1681620392
transform 1 0 2660 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1852
timestamp 1681620392
transform 1 0 2692 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_2154
timestamp 1681620392
transform 1 0 2692 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1817
timestamp 1681620392
transform 1 0 2708 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_2245
timestamp 1681620392
transform 1 0 2700 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2246
timestamp 1681620392
transform 1 0 2708 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2247
timestamp 1681620392
transform 1 0 2716 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2337
timestamp 1681620392
transform 1 0 2700 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1949
timestamp 1681620392
transform 1 0 2700 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_2248
timestamp 1681620392
transform 1 0 2740 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2338
timestamp 1681620392
transform 1 0 2732 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2155
timestamp 1681620392
transform 1 0 2748 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1880
timestamp 1681620392
transform 1 0 2764 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1824
timestamp 1681620392
transform 1 0 2812 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_2126
timestamp 1681620392
transform 1 0 2788 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_2156
timestamp 1681620392
transform 1 0 2780 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2157
timestamp 1681620392
transform 1 0 2796 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_1906
timestamp 1681620392
transform 1 0 2748 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_2249
timestamp 1681620392
transform 1 0 2764 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2250
timestamp 1681620392
transform 1 0 2772 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1907
timestamp 1681620392
transform 1 0 2780 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1881
timestamp 1681620392
transform 1 0 2812 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1825
timestamp 1681620392
transform 1 0 2860 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1853
timestamp 1681620392
transform 1 0 2852 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_2158
timestamp 1681620392
transform 1 0 2836 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2251
timestamp 1681620392
transform 1 0 2796 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2252
timestamp 1681620392
transform 1 0 2812 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2253
timestamp 1681620392
transform 1 0 2820 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_1969
timestamp 1681620392
transform 1 0 2804 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_2254
timestamp 1681620392
transform 1 0 2844 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2255
timestamp 1681620392
transform 1 0 2852 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2256
timestamp 1681620392
transform 1 0 2868 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2339
timestamp 1681620392
transform 1 0 2836 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2340
timestamp 1681620392
transform 1 0 2844 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1950
timestamp 1681620392
transform 1 0 2836 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_2341
timestamp 1681620392
transform 1 0 2876 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_1951
timestamp 1681620392
transform 1 0 2876 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1970
timestamp 1681620392
transform 1 0 2876 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1854
timestamp 1681620392
transform 1 0 2916 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_2159
timestamp 1681620392
transform 1 0 2916 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2342
timestamp 1681620392
transform 1 0 2916 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2160
timestamp 1681620392
transform 1 0 2948 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2343
timestamp 1681620392
transform 1 0 2956 0 1 1805
box -2 -2 2 2
use Project_Top_VIA0  Project_Top_VIA0_24
timestamp 1681620392
transform 1 0 48 0 1 1770
box -10 -3 10 3
use FILL  FILL_463
timestamp 1681620392
transform 1 0 72 0 1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_144
timestamp 1681620392
transform 1 0 80 0 1 1770
box -8 -3 34 105
use INVX2  INVX2_138
timestamp 1681620392
transform -1 0 128 0 1 1770
box -9 -3 26 105
use FILL  FILL_464
timestamp 1681620392
transform 1 0 128 0 1 1770
box -8 -3 16 105
use FILL  FILL_465
timestamp 1681620392
transform 1 0 136 0 1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_145
timestamp 1681620392
transform 1 0 144 0 1 1770
box -8 -3 34 105
use NOR2X1  NOR2X1_39
timestamp 1681620392
transform 1 0 176 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_40
timestamp 1681620392
transform -1 0 224 0 1 1770
box -8 -3 32 105
use INVX2  INVX2_139
timestamp 1681620392
transform 1 0 224 0 1 1770
box -9 -3 26 105
use FILL  FILL_466
timestamp 1681620392
transform 1 0 240 0 1 1770
box -8 -3 16 105
use FILL  FILL_467
timestamp 1681620392
transform 1 0 248 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_140
timestamp 1681620392
transform -1 0 272 0 1 1770
box -9 -3 26 105
use NAND2X1  NAND2X1_120
timestamp 1681620392
transform 1 0 272 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_121
timestamp 1681620392
transform 1 0 296 0 1 1770
box -8 -3 32 105
use OAI21X1  OAI21X1_146
timestamp 1681620392
transform -1 0 352 0 1 1770
box -8 -3 34 105
use NAND2X1  NAND2X1_122
timestamp 1681620392
transform 1 0 352 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_123
timestamp 1681620392
transform 1 0 376 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_124
timestamp 1681620392
transform 1 0 400 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_125
timestamp 1681620392
transform -1 0 448 0 1 1770
box -8 -3 32 105
use OAI21X1  OAI21X1_147
timestamp 1681620392
transform 1 0 448 0 1 1770
box -8 -3 34 105
use NAND2X1  NAND2X1_126
timestamp 1681620392
transform 1 0 480 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_41
timestamp 1681620392
transform 1 0 504 0 1 1770
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_140
timestamp 1681620392
transform 1 0 528 0 1 1770
box -8 -3 104 105
use OAI22X1  OAI22X1_22
timestamp 1681620392
transform -1 0 664 0 1 1770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_141
timestamp 1681620392
transform 1 0 664 0 1 1770
box -8 -3 104 105
use INVX2  INVX2_142
timestamp 1681620392
transform 1 0 760 0 1 1770
box -9 -3 26 105
use M3_M2  M3_M2_1971
timestamp 1681620392
transform 1 0 796 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1972
timestamp 1681620392
transform 1 0 820 0 1 1775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_142
timestamp 1681620392
transform 1 0 776 0 1 1770
box -8 -3 104 105
use NAND2X1  NAND2X1_127
timestamp 1681620392
transform -1 0 896 0 1 1770
box -8 -3 32 105
use NAND3X1  NAND3X1_48
timestamp 1681620392
transform -1 0 928 0 1 1770
box -8 -3 40 105
use AND2X2  AND2X2_12
timestamp 1681620392
transform 1 0 928 0 1 1770
box -8 -3 40 105
use INVX2  INVX2_143
timestamp 1681620392
transform -1 0 976 0 1 1770
box -9 -3 26 105
use OAI22X1  OAI22X1_23
timestamp 1681620392
transform -1 0 1016 0 1 1770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_143
timestamp 1681620392
transform -1 0 1112 0 1 1770
box -8 -3 104 105
use NAND3X1  NAND3X1_49
timestamp 1681620392
transform 1 0 1112 0 1 1770
box -8 -3 40 105
use INVX2  INVX2_144
timestamp 1681620392
transform 1 0 1144 0 1 1770
box -9 -3 26 105
use M3_M2  M3_M2_1973
timestamp 1681620392
transform 1 0 1196 0 1 1775
box -3 -3 3 3
use NAND3X1  NAND3X1_50
timestamp 1681620392
transform 1 0 1160 0 1 1770
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_144
timestamp 1681620392
transform 1 0 1192 0 1 1770
box -8 -3 104 105
use M3_M2  M3_M2_1974
timestamp 1681620392
transform 1 0 1316 0 1 1775
box -3 -3 3 3
use NAND2X1  NAND2X1_128
timestamp 1681620392
transform 1 0 1288 0 1 1770
box -8 -3 32 105
use AND2X2  AND2X2_13
timestamp 1681620392
transform -1 0 1344 0 1 1770
box -8 -3 40 105
use M3_M2  M3_M2_1975
timestamp 1681620392
transform 1 0 1372 0 1 1775
box -3 -3 3 3
use NOR2X1  NOR2X1_42
timestamp 1681620392
transform -1 0 1368 0 1 1770
box -8 -3 32 105
use FILL  FILL_477
timestamp 1681620392
transform 1 0 1368 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_145
timestamp 1681620392
transform 1 0 1376 0 1 1770
box -9 -3 26 105
use FILL  FILL_478
timestamp 1681620392
transform 1 0 1392 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_16
timestamp 1681620392
transform 1 0 1400 0 1 1770
box -5 -3 28 105
use OAI21X1  OAI21X1_152
timestamp 1681620392
transform 1 0 1424 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_153
timestamp 1681620392
transform 1 0 1456 0 1 1770
box -8 -3 34 105
use OAI22X1  OAI22X1_24
timestamp 1681620392
transform -1 0 1528 0 1 1770
box -8 -3 46 105
use INVX2  INVX2_146
timestamp 1681620392
transform -1 0 1544 0 1 1770
box -9 -3 26 105
use NAND2X1  NAND2X1_129
timestamp 1681620392
transform -1 0 1568 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_130
timestamp 1681620392
transform 1 0 1568 0 1 1770
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_145
timestamp 1681620392
transform -1 0 1688 0 1 1770
box -8 -3 104 105
use OAI21X1  OAI21X1_154
timestamp 1681620392
transform 1 0 1688 0 1 1770
box -8 -3 34 105
use FILL  FILL_479
timestamp 1681620392
transform 1 0 1720 0 1 1770
box -8 -3 16 105
use FILL  FILL_505
timestamp 1681620392
transform 1 0 1728 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_1976
timestamp 1681620392
transform 1 0 1772 0 1 1775
box -3 -3 3 3
use OAI22X1  OAI22X1_30
timestamp 1681620392
transform 1 0 1736 0 1 1770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_148
timestamp 1681620392
transform 1 0 1776 0 1 1770
box -8 -3 104 105
use INVX2  INVX2_157
timestamp 1681620392
transform 1 0 1872 0 1 1770
box -9 -3 26 105
use M3_M2  M3_M2_1977
timestamp 1681620392
transform 1 0 1908 0 1 1775
box -3 -3 3 3
use NAND2X1  NAND2X1_138
timestamp 1681620392
transform 1 0 1888 0 1 1770
box -8 -3 32 105
use FILL  FILL_507
timestamp 1681620392
transform 1 0 1912 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_31
timestamp 1681620392
transform -1 0 1960 0 1 1770
box -8 -3 46 105
use INVX2  INVX2_158
timestamp 1681620392
transform -1 0 1976 0 1 1770
box -9 -3 26 105
use FILL  FILL_508
timestamp 1681620392
transform 1 0 1976 0 1 1770
box -8 -3 16 105
use FILL  FILL_509
timestamp 1681620392
transform 1 0 1984 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_1978
timestamp 1681620392
transform 1 0 2020 0 1 1775
box -3 -3 3 3
use OAI22X1  OAI22X1_32
timestamp 1681620392
transform -1 0 2032 0 1 1770
box -8 -3 46 105
use M3_M2  M3_M2_1979
timestamp 1681620392
transform 1 0 2044 0 1 1775
box -3 -3 3 3
use FILL  FILL_510
timestamp 1681620392
transform 1 0 2032 0 1 1770
box -8 -3 16 105
use NAND2X1  NAND2X1_139
timestamp 1681620392
transform 1 0 2040 0 1 1770
box -8 -3 32 105
use INVX2  INVX2_159
timestamp 1681620392
transform -1 0 2080 0 1 1770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_149
timestamp 1681620392
transform 1 0 2080 0 1 1770
box -8 -3 104 105
use INVX2  INVX2_160
timestamp 1681620392
transform 1 0 2176 0 1 1770
box -9 -3 26 105
use FILL  FILL_511
timestamp 1681620392
transform 1 0 2192 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_150
timestamp 1681620392
transform 1 0 2200 0 1 1770
box -8 -3 104 105
use OAI22X1  OAI22X1_33
timestamp 1681620392
transform -1 0 2336 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_34
timestamp 1681620392
transform -1 0 2376 0 1 1770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_151
timestamp 1681620392
transform 1 0 2376 0 1 1770
box -8 -3 104 105
use INVX2  INVX2_161
timestamp 1681620392
transform 1 0 2472 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_162
timestamp 1681620392
transform 1 0 2488 0 1 1770
box -9 -3 26 105
use OAI21X1  OAI21X1_157
timestamp 1681620392
transform 1 0 2504 0 1 1770
box -8 -3 34 105
use FILL  FILL_512
timestamp 1681620392
transform 1 0 2536 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_17
timestamp 1681620392
transform -1 0 2568 0 1 1770
box -5 -3 28 105
use FILL  FILL_513
timestamp 1681620392
transform 1 0 2568 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_163
timestamp 1681620392
transform -1 0 2592 0 1 1770
box -9 -3 26 105
use FILL  FILL_514
timestamp 1681620392
transform 1 0 2592 0 1 1770
box -8 -3 16 105
use FILL  FILL_515
timestamp 1681620392
transform 1 0 2600 0 1 1770
box -8 -3 16 105
use NAND2X1  NAND2X1_140
timestamp 1681620392
transform -1 0 2632 0 1 1770
box -8 -3 32 105
use AOI21X1  AOI21X1_12
timestamp 1681620392
transform -1 0 2664 0 1 1770
box -7 -3 39 105
use OAI21X1  OAI21X1_158
timestamp 1681620392
transform 1 0 2664 0 1 1770
box -8 -3 34 105
use INVX2  INVX2_164
timestamp 1681620392
transform 1 0 2696 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_165
timestamp 1681620392
transform 1 0 2712 0 1 1770
box -9 -3 26 105
use FILL  FILL_516
timestamp 1681620392
transform 1 0 2728 0 1 1770
box -8 -3 16 105
use FILL  FILL_517
timestamp 1681620392
transform 1 0 2736 0 1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_159
timestamp 1681620392
transform -1 0 2776 0 1 1770
box -8 -3 34 105
use NAND3X1  NAND3X1_52
timestamp 1681620392
transform -1 0 2808 0 1 1770
box -8 -3 40 105
use OAI21X1  OAI21X1_160
timestamp 1681620392
transform 1 0 2808 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_161
timestamp 1681620392
transform 1 0 2840 0 1 1770
box -8 -3 34 105
use FILL  FILL_518
timestamp 1681620392
transform 1 0 2872 0 1 1770
box -8 -3 16 105
use FILL  FILL_519
timestamp 1681620392
transform 1 0 2880 0 1 1770
box -8 -3 16 105
use FILL  FILL_520
timestamp 1681620392
transform 1 0 2888 0 1 1770
box -8 -3 16 105
use NAND2X1  NAND2X1_141
timestamp 1681620392
transform 1 0 2896 0 1 1770
box -8 -3 32 105
use OAI21X1  OAI21X1_162
timestamp 1681620392
transform 1 0 2920 0 1 1770
box -8 -3 34 105
use FILL  FILL_521
timestamp 1681620392
transform 1 0 2952 0 1 1770
box -8 -3 16 105
use FILL  FILL_522
timestamp 1681620392
transform 1 0 2960 0 1 1770
box -8 -3 16 105
use FILL  FILL_523
timestamp 1681620392
transform 1 0 2968 0 1 1770
box -8 -3 16 105
use FILL  FILL_524
timestamp 1681620392
transform 1 0 2976 0 1 1770
box -8 -3 16 105
use FILL  FILL_525
timestamp 1681620392
transform 1 0 2984 0 1 1770
box -8 -3 16 105
use FILL  FILL_526
timestamp 1681620392
transform 1 0 2992 0 1 1770
box -8 -3 16 105
use FILL  FILL_527
timestamp 1681620392
transform 1 0 3000 0 1 1770
box -8 -3 16 105
use FILL  FILL_528
timestamp 1681620392
transform 1 0 3008 0 1 1770
box -8 -3 16 105
use Project_Top_VIA0  Project_Top_VIA0_25
timestamp 1681620392
transform 1 0 3043 0 1 1770
box -10 -3 10 3
use M3_M2  M3_M2_1980
timestamp 1681620392
transform 1 0 84 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1998
timestamp 1681620392
transform 1 0 76 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1999
timestamp 1681620392
transform 1 0 124 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2014
timestamp 1681620392
transform 1 0 116 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2358
timestamp 1681620392
transform 1 0 84 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_2044
timestamp 1681620392
transform 1 0 172 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_2359
timestamp 1681620392
transform 1 0 180 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2437
timestamp 1681620392
transform 1 0 108 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2438
timestamp 1681620392
transform 1 0 164 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2096
timestamp 1681620392
transform 1 0 68 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1981
timestamp 1681620392
transform 1 0 196 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_2439
timestamp 1681620392
transform 1 0 204 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2097
timestamp 1681620392
transform 1 0 204 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1982
timestamp 1681620392
transform 1 0 228 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2000
timestamp 1681620392
transform 1 0 220 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_2360
timestamp 1681620392
transform 1 0 220 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_2045
timestamp 1681620392
transform 1 0 244 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2046
timestamp 1681620392
transform 1 0 268 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2047
timestamp 1681620392
transform 1 0 300 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2066
timestamp 1681620392
transform 1 0 220 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_2440
timestamp 1681620392
transform 1 0 244 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2067
timestamp 1681620392
transform 1 0 260 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2015
timestamp 1681620392
transform 1 0 316 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2361
timestamp 1681620392
transform 1 0 316 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2441
timestamp 1681620392
transform 1 0 300 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2068
timestamp 1681620392
transform 1 0 308 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2098
timestamp 1681620392
transform 1 0 308 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2069
timestamp 1681620392
transform 1 0 324 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_2362
timestamp 1681620392
transform 1 0 348 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2363
timestamp 1681620392
transform 1 0 364 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2442
timestamp 1681620392
transform 1 0 340 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2522
timestamp 1681620392
transform 1 0 324 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_2070
timestamp 1681620392
transform 1 0 356 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_2523
timestamp 1681620392
transform 1 0 356 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_2118
timestamp 1681620392
transform 1 0 356 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_2364
timestamp 1681620392
transform 1 0 396 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2365
timestamp 1681620392
transform 1 0 420 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2443
timestamp 1681620392
transform 1 0 380 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2444
timestamp 1681620392
transform 1 0 396 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2445
timestamp 1681620392
transform 1 0 412 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2524
timestamp 1681620392
transform 1 0 396 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_2119
timestamp 1681620392
transform 1 0 396 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_2446
timestamp 1681620392
transform 1 0 436 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2366
timestamp 1681620392
transform 1 0 452 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_2048
timestamp 1681620392
transform 1 0 468 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2016
timestamp 1681620392
transform 1 0 492 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2017
timestamp 1681620392
transform 1 0 524 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2367
timestamp 1681620392
transform 1 0 476 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2368
timestamp 1681620392
transform 1 0 484 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2369
timestamp 1681620392
transform 1 0 500 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2370
timestamp 1681620392
transform 1 0 516 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2371
timestamp 1681620392
transform 1 0 524 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_2071
timestamp 1681620392
transform 1 0 484 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_2447
timestamp 1681620392
transform 1 0 492 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2448
timestamp 1681620392
transform 1 0 508 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2449
timestamp 1681620392
transform 1 0 524 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2525
timestamp 1681620392
transform 1 0 476 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_2099
timestamp 1681620392
transform 1 0 508 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2120
timestamp 1681620392
transform 1 0 476 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2140
timestamp 1681620392
transform 1 0 508 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2001
timestamp 1681620392
transform 1 0 540 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_2450
timestamp 1681620392
transform 1 0 548 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2002
timestamp 1681620392
transform 1 0 564 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2018
timestamp 1681620392
transform 1 0 588 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2372
timestamp 1681620392
transform 1 0 564 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2373
timestamp 1681620392
transform 1 0 580 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2451
timestamp 1681620392
transform 1 0 572 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2452
timestamp 1681620392
transform 1 0 588 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2148
timestamp 1681620392
transform 1 0 572 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2003
timestamp 1681620392
transform 1 0 628 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2019
timestamp 1681620392
transform 1 0 620 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2374
timestamp 1681620392
transform 1 0 620 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1983
timestamp 1681620392
transform 1 0 636 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_2349
timestamp 1681620392
transform 1 0 660 0 1 1745
box -2 -2 2 2
use M3_M2  M3_M2_2072
timestamp 1681620392
transform 1 0 652 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_2350
timestamp 1681620392
transform 1 0 684 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_2453
timestamp 1681620392
transform 1 0 684 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2100
timestamp 1681620392
transform 1 0 684 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_2351
timestamp 1681620392
transform 1 0 700 0 1 1745
box -2 -2 2 2
use M3_M2  M3_M2_2020
timestamp 1681620392
transform 1 0 708 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2375
timestamp 1681620392
transform 1 0 700 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2454
timestamp 1681620392
transform 1 0 708 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2121
timestamp 1681620392
transform 1 0 708 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_2352
timestamp 1681620392
transform 1 0 724 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_2376
timestamp 1681620392
transform 1 0 732 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2377
timestamp 1681620392
transform 1 0 740 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2455
timestamp 1681620392
transform 1 0 724 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2073
timestamp 1681620392
transform 1 0 732 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2101
timestamp 1681620392
transform 1 0 724 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2122
timestamp 1681620392
transform 1 0 740 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_2353
timestamp 1681620392
transform 1 0 764 0 1 1745
box -2 -2 2 2
use M3_M2  M3_M2_2021
timestamp 1681620392
transform 1 0 780 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2378
timestamp 1681620392
transform 1 0 772 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2456
timestamp 1681620392
transform 1 0 764 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2022
timestamp 1681620392
transform 1 0 820 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2379
timestamp 1681620392
transform 1 0 796 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2380
timestamp 1681620392
transform 1 0 804 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_2049
timestamp 1681620392
transform 1 0 812 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_2457
timestamp 1681620392
transform 1 0 780 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2458
timestamp 1681620392
transform 1 0 788 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2074
timestamp 1681620392
transform 1 0 804 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2123
timestamp 1681620392
transform 1 0 772 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2023
timestamp 1681620392
transform 1 0 844 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2381
timestamp 1681620392
transform 1 0 844 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2382
timestamp 1681620392
transform 1 0 852 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2459
timestamp 1681620392
transform 1 0 820 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2460
timestamp 1681620392
transform 1 0 836 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2075
timestamp 1681620392
transform 1 0 844 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_2526
timestamp 1681620392
transform 1 0 820 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_2102
timestamp 1681620392
transform 1 0 836 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_2527
timestamp 1681620392
transform 1 0 844 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_2124
timestamp 1681620392
transform 1 0 844 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2004
timestamp 1681620392
transform 1 0 876 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_2354
timestamp 1681620392
transform 1 0 868 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_2383
timestamp 1681620392
transform 1 0 884 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2384
timestamp 1681620392
transform 1 0 892 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2461
timestamp 1681620392
transform 1 0 860 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2462
timestamp 1681620392
transform 1 0 868 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2076
timestamp 1681620392
transform 1 0 884 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2103
timestamp 1681620392
transform 1 0 876 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2005
timestamp 1681620392
transform 1 0 924 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2024
timestamp 1681620392
transform 1 0 972 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2385
timestamp 1681620392
transform 1 0 932 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2386
timestamp 1681620392
transform 1 0 1020 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2463
timestamp 1681620392
transform 1 0 908 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2077
timestamp 1681620392
transform 1 0 916 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2050
timestamp 1681620392
transform 1 0 1028 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1984
timestamp 1681620392
transform 1 0 1068 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2025
timestamp 1681620392
transform 1 0 1076 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2387
timestamp 1681620392
transform 1 0 1036 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2388
timestamp 1681620392
transform 1 0 1052 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2389
timestamp 1681620392
transform 1 0 1076 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2464
timestamp 1681620392
transform 1 0 972 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2465
timestamp 1681620392
transform 1 0 1020 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2466
timestamp 1681620392
transform 1 0 1028 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2467
timestamp 1681620392
transform 1 0 1044 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2528
timestamp 1681620392
transform 1 0 916 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_2125
timestamp 1681620392
transform 1 0 916 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2104
timestamp 1681620392
transform 1 0 1020 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2141
timestamp 1681620392
transform 1 0 1044 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2051
timestamp 1681620392
transform 1 0 1084 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_2390
timestamp 1681620392
transform 1 0 1092 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2468
timestamp 1681620392
transform 1 0 1068 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2469
timestamp 1681620392
transform 1 0 1084 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2126
timestamp 1681620392
transform 1 0 1092 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_2391
timestamp 1681620392
transform 1 0 1116 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2392
timestamp 1681620392
transform 1 0 1132 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_2052
timestamp 1681620392
transform 1 0 1140 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_2393
timestamp 1681620392
transform 1 0 1148 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2394
timestamp 1681620392
transform 1 0 1156 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2470
timestamp 1681620392
transform 1 0 1108 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2471
timestamp 1681620392
transform 1 0 1124 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2472
timestamp 1681620392
transform 1 0 1140 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2473
timestamp 1681620392
transform 1 0 1148 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2078
timestamp 1681620392
transform 1 0 1156 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2127
timestamp 1681620392
transform 1 0 1148 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2149
timestamp 1681620392
transform 1 0 1124 0 1 1685
box -3 -3 3 3
use M2_M1  M2_M1_2355
timestamp 1681620392
transform 1 0 1172 0 1 1745
box -2 -2 2 2
use M3_M2  M3_M2_2053
timestamp 1681620392
transform 1 0 1172 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_2395
timestamp 1681620392
transform 1 0 1196 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_2054
timestamp 1681620392
transform 1 0 1204 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_2396
timestamp 1681620392
transform 1 0 1212 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_2079
timestamp 1681620392
transform 1 0 1188 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_2474
timestamp 1681620392
transform 1 0 1196 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2475
timestamp 1681620392
transform 1 0 1204 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2105
timestamp 1681620392
transform 1 0 1212 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2142
timestamp 1681620392
transform 1 0 1188 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_2356
timestamp 1681620392
transform 1 0 1236 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_2397
timestamp 1681620392
transform 1 0 1244 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_2128
timestamp 1681620392
transform 1 0 1236 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1985
timestamp 1681620392
transform 1 0 1276 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1986
timestamp 1681620392
transform 1 0 1292 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2006
timestamp 1681620392
transform 1 0 1268 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2026
timestamp 1681620392
transform 1 0 1260 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2476
timestamp 1681620392
transform 1 0 1260 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2106
timestamp 1681620392
transform 1 0 1260 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2150
timestamp 1681620392
transform 1 0 1252 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2027
timestamp 1681620392
transform 1 0 1284 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2357
timestamp 1681620392
transform 1 0 1300 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_2398
timestamp 1681620392
transform 1 0 1284 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2477
timestamp 1681620392
transform 1 0 1276 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2080
timestamp 1681620392
transform 1 0 1284 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_2478
timestamp 1681620392
transform 1 0 1300 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2479
timestamp 1681620392
transform 1 0 1308 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2143
timestamp 1681620392
transform 1 0 1276 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2107
timestamp 1681620392
transform 1 0 1300 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2129
timestamp 1681620392
transform 1 0 1308 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2007
timestamp 1681620392
transform 1 0 1324 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_2399
timestamp 1681620392
transform 1 0 1316 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2400
timestamp 1681620392
transform 1 0 1324 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2480
timestamp 1681620392
transform 1 0 1324 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2081
timestamp 1681620392
transform 1 0 1332 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_2481
timestamp 1681620392
transform 1 0 1340 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2130
timestamp 1681620392
transform 1 0 1324 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_2529
timestamp 1681620392
transform 1 0 1340 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_2108
timestamp 1681620392
transform 1 0 1348 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_2544
timestamp 1681620392
transform 1 0 1348 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_2055
timestamp 1681620392
transform 1 0 1396 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_2401
timestamp 1681620392
transform 1 0 1404 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2402
timestamp 1681620392
transform 1 0 1412 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2482
timestamp 1681620392
transform 1 0 1364 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2082
timestamp 1681620392
transform 1 0 1380 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_2530
timestamp 1681620392
transform 1 0 1380 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2531
timestamp 1681620392
transform 1 0 1388 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_2131
timestamp 1681620392
transform 1 0 1364 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_2483
timestamp 1681620392
transform 1 0 1404 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2083
timestamp 1681620392
transform 1 0 1412 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_2484
timestamp 1681620392
transform 1 0 1452 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2008
timestamp 1681620392
transform 1 0 1468 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2009
timestamp 1681620392
transform 1 0 1508 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1987
timestamp 1681620392
transform 1 0 1572 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_2403
timestamp 1681620392
transform 1 0 1476 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2404
timestamp 1681620392
transform 1 0 1564 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2485
timestamp 1681620392
transform 1 0 1500 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2486
timestamp 1681620392
transform 1 0 1556 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2487
timestamp 1681620392
transform 1 0 1580 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2532
timestamp 1681620392
transform 1 0 1564 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_2132
timestamp 1681620392
transform 1 0 1564 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2151
timestamp 1681620392
transform 1 0 1532 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2084
timestamp 1681620392
transform 1 0 1588 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_2405
timestamp 1681620392
transform 1 0 1620 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1988
timestamp 1681620392
transform 1 0 1652 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_2406
timestamp 1681620392
transform 1 0 1636 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_2085
timestamp 1681620392
transform 1 0 1636 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_2488
timestamp 1681620392
transform 1 0 1644 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2533
timestamp 1681620392
transform 1 0 1636 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_2109
timestamp 1681620392
transform 1 0 1644 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1989
timestamp 1681620392
transform 1 0 1668 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2028
timestamp 1681620392
transform 1 0 1660 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2407
timestamp 1681620392
transform 1 0 1668 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2489
timestamp 1681620392
transform 1 0 1660 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2490
timestamp 1681620392
transform 1 0 1668 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2534
timestamp 1681620392
transform 1 0 1660 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_2110
timestamp 1681620392
transform 1 0 1668 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2029
timestamp 1681620392
transform 1 0 1700 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2086
timestamp 1681620392
transform 1 0 1692 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_2535
timestamp 1681620392
transform 1 0 1700 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_2111
timestamp 1681620392
transform 1 0 1708 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2133
timestamp 1681620392
transform 1 0 1700 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2056
timestamp 1681620392
transform 1 0 1724 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_2536
timestamp 1681620392
transform 1 0 1732 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_2010
timestamp 1681620392
transform 1 0 1748 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2011
timestamp 1681620392
transform 1 0 1780 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_2408
timestamp 1681620392
transform 1 0 1740 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2409
timestamp 1681620392
transform 1 0 1748 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2410
timestamp 1681620392
transform 1 0 1764 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_2057
timestamp 1681620392
transform 1 0 1772 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_2411
timestamp 1681620392
transform 1 0 1796 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2491
timestamp 1681620392
transform 1 0 1756 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2492
timestamp 1681620392
transform 1 0 1772 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2412
timestamp 1681620392
transform 1 0 1836 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1990
timestamp 1681620392
transform 1 0 1860 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2030
timestamp 1681620392
transform 1 0 1868 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2413
timestamp 1681620392
transform 1 0 1868 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2493
timestamp 1681620392
transform 1 0 1844 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2494
timestamp 1681620392
transform 1 0 1860 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2495
timestamp 1681620392
transform 1 0 1868 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2537
timestamp 1681620392
transform 1 0 1844 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2538
timestamp 1681620392
transform 1 0 1876 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1991
timestamp 1681620392
transform 1 0 1932 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2012
timestamp 1681620392
transform 1 0 1996 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2031
timestamp 1681620392
transform 1 0 1908 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2414
timestamp 1681620392
transform 1 0 1892 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2415
timestamp 1681620392
transform 1 0 1908 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_2087
timestamp 1681620392
transform 1 0 1908 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1992
timestamp 1681620392
transform 1 0 2100 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2032
timestamp 1681620392
transform 1 0 2004 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2033
timestamp 1681620392
transform 1 0 2092 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2416
timestamp 1681620392
transform 1 0 2004 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2417
timestamp 1681620392
transform 1 0 2092 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2496
timestamp 1681620392
transform 1 0 1940 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2497
timestamp 1681620392
transform 1 0 1988 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2498
timestamp 1681620392
transform 1 0 2028 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2088
timestamp 1681620392
transform 1 0 2052 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_2499
timestamp 1681620392
transform 1 0 2084 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2089
timestamp 1681620392
transform 1 0 2092 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2112
timestamp 1681620392
transform 1 0 1988 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2134
timestamp 1681620392
transform 1 0 1900 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2135
timestamp 1681620392
transform 1 0 1956 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2144
timestamp 1681620392
transform 1 0 1884 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2152
timestamp 1681620392
transform 1 0 1876 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2145
timestamp 1681620392
transform 1 0 1924 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2153
timestamp 1681620392
transform 1 0 1908 0 1 1685
box -3 -3 3 3
use M2_M1  M2_M1_2539
timestamp 1681620392
transform 1 0 2108 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1993
timestamp 1681620392
transform 1 0 2124 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_2500
timestamp 1681620392
transform 1 0 2124 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2034
timestamp 1681620392
transform 1 0 2172 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2035
timestamp 1681620392
transform 1 0 2212 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2418
timestamp 1681620392
transform 1 0 2172 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_2058
timestamp 1681620392
transform 1 0 2196 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2090
timestamp 1681620392
transform 1 0 2172 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_2501
timestamp 1681620392
transform 1 0 2196 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2091
timestamp 1681620392
transform 1 0 2260 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2113
timestamp 1681620392
transform 1 0 2252 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_2502
timestamp 1681620392
transform 1 0 2276 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2419
timestamp 1681620392
transform 1 0 2284 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_2013
timestamp 1681620392
transform 1 0 2300 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2036
timestamp 1681620392
transform 1 0 2332 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2420
timestamp 1681620392
transform 1 0 2324 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2421
timestamp 1681620392
transform 1 0 2340 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2503
timestamp 1681620392
transform 1 0 2316 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2059
timestamp 1681620392
transform 1 0 2356 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_2504
timestamp 1681620392
transform 1 0 2348 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2092
timestamp 1681620392
transform 1 0 2356 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_2422
timestamp 1681620392
transform 1 0 2372 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1994
timestamp 1681620392
transform 1 0 2388 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2037
timestamp 1681620392
transform 1 0 2460 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2423
timestamp 1681620392
transform 1 0 2388 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_2060
timestamp 1681620392
transform 1 0 2412 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2061
timestamp 1681620392
transform 1 0 2468 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_2424
timestamp 1681620392
transform 1 0 2484 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2505
timestamp 1681620392
transform 1 0 2412 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2506
timestamp 1681620392
transform 1 0 2468 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2507
timestamp 1681620392
transform 1 0 2476 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2154
timestamp 1681620392
transform 1 0 2428 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2155
timestamp 1681620392
transform 1 0 2444 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2062
timestamp 1681620392
transform 1 0 2492 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2114
timestamp 1681620392
transform 1 0 2492 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1995
timestamp 1681620392
transform 1 0 2556 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2038
timestamp 1681620392
transform 1 0 2556 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2039
timestamp 1681620392
transform 1 0 2596 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2425
timestamp 1681620392
transform 1 0 2508 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2426
timestamp 1681620392
transform 1 0 2596 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2508
timestamp 1681620392
transform 1 0 2556 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2509
timestamp 1681620392
transform 1 0 2588 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2427
timestamp 1681620392
transform 1 0 2620 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2428
timestamp 1681620392
transform 1 0 2628 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2510
timestamp 1681620392
transform 1 0 2612 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2511
timestamp 1681620392
transform 1 0 2620 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2115
timestamp 1681620392
transform 1 0 2588 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_2540
timestamp 1681620392
transform 1 0 2596 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_2156
timestamp 1681620392
transform 1 0 2508 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2157
timestamp 1681620392
transform 1 0 2564 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2116
timestamp 1681620392
transform 1 0 2628 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2136
timestamp 1681620392
transform 1 0 2612 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2137
timestamp 1681620392
transform 1 0 2628 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_2429
timestamp 1681620392
transform 1 0 2740 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2512
timestamp 1681620392
transform 1 0 2660 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2513
timestamp 1681620392
transform 1 0 2716 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2430
timestamp 1681620392
transform 1 0 2756 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_1996
timestamp 1681620392
transform 1 0 2772 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2040
timestamp 1681620392
transform 1 0 2788 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2431
timestamp 1681620392
transform 1 0 2788 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2432
timestamp 1681620392
transform 1 0 2796 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2514
timestamp 1681620392
transform 1 0 2772 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2541
timestamp 1681620392
transform 1 0 2788 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_1997
timestamp 1681620392
transform 1 0 2820 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2041
timestamp 1681620392
transform 1 0 2812 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2433
timestamp 1681620392
transform 1 0 2812 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2515
timestamp 1681620392
transform 1 0 2812 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2042
timestamp 1681620392
transform 1 0 2868 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2434
timestamp 1681620392
transform 1 0 2876 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_2093
timestamp 1681620392
transform 1 0 2860 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2043
timestamp 1681620392
transform 1 0 2948 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_2435
timestamp 1681620392
transform 1 0 2908 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2516
timestamp 1681620392
transform 1 0 2868 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2517
timestamp 1681620392
transform 1 0 2876 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_2094
timestamp 1681620392
transform 1 0 2884 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2095
timestamp 1681620392
transform 1 0 2900 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2063
timestamp 1681620392
transform 1 0 2916 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_2436
timestamp 1681620392
transform 1 0 2932 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_2064
timestamp 1681620392
transform 1 0 2972 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2065
timestamp 1681620392
transform 1 0 3012 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_2518
timestamp 1681620392
transform 1 0 2908 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2519
timestamp 1681620392
transform 1 0 2916 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2520
timestamp 1681620392
transform 1 0 2956 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2521
timestamp 1681620392
transform 1 0 3012 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2542
timestamp 1681620392
transform 1 0 2868 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_2138
timestamp 1681620392
transform 1 0 2860 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_2543
timestamp 1681620392
transform 1 0 2900 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_2139
timestamp 1681620392
transform 1 0 2900 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2117
timestamp 1681620392
transform 1 0 2916 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2146
timestamp 1681620392
transform 1 0 2908 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2147
timestamp 1681620392
transform 1 0 2956 0 1 1695
box -3 -3 3 3
use Project_Top_VIA0  Project_Top_VIA0_26
timestamp 1681620392
transform 1 0 24 0 1 1670
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_138
timestamp 1681620392
transform 1 0 72 0 -1 1770
box -8 -3 104 105
use FILL  FILL_468
timestamp 1681620392
transform 1 0 168 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_141
timestamp 1681620392
transform 1 0 176 0 -1 1770
box -9 -3 26 105
use FILL  FILL_469
timestamp 1681620392
transform 1 0 192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_470
timestamp 1681620392
transform 1 0 200 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_139
timestamp 1681620392
transform 1 0 208 0 -1 1770
box -8 -3 104 105
use FILL  FILL_471
timestamp 1681620392
transform 1 0 304 0 -1 1770
box -8 -3 16 105
use FILL  FILL_472
timestamp 1681620392
transform 1 0 312 0 -1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_148
timestamp 1681620392
transform -1 0 352 0 -1 1770
box -8 -3 34 105
use FILL  FILL_473
timestamp 1681620392
transform 1 0 352 0 -1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_149
timestamp 1681620392
transform -1 0 392 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_150
timestamp 1681620392
transform -1 0 424 0 -1 1770
box -8 -3 34 105
use FILL  FILL_474
timestamp 1681620392
transform 1 0 424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_475
timestamp 1681620392
transform 1 0 432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_476
timestamp 1681620392
transform 1 0 440 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_2158
timestamp 1681620392
transform 1 0 460 0 1 1675
box -3 -3 3 3
use OAI21X1  OAI21X1_151
timestamp 1681620392
transform 1 0 448 0 -1 1770
box -8 -3 34 105
use OAI22X1  OAI22X1_25
timestamp 1681620392
transform 1 0 480 0 -1 1770
box -8 -3 46 105
use INVX2  INVX2_147
timestamp 1681620392
transform 1 0 520 0 -1 1770
box -9 -3 26 105
use FILL  FILL_480
timestamp 1681620392
transform 1 0 536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_481
timestamp 1681620392
transform 1 0 544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_482
timestamp 1681620392
transform 1 0 552 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_26
timestamp 1681620392
transform -1 0 600 0 -1 1770
box -8 -3 46 105
use FILL  FILL_483
timestamp 1681620392
transform 1 0 600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_484
timestamp 1681620392
transform 1 0 608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_485
timestamp 1681620392
transform 1 0 616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_486
timestamp 1681620392
transform 1 0 624 0 -1 1770
box -8 -3 16 105
use FILL  FILL_487
timestamp 1681620392
transform 1 0 632 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_148
timestamp 1681620392
transform 1 0 640 0 -1 1770
box -9 -3 26 105
use FILL  FILL_488
timestamp 1681620392
transform 1 0 656 0 -1 1770
box -8 -3 16 105
use FILL  FILL_489
timestamp 1681620392
transform 1 0 664 0 -1 1770
box -8 -3 16 105
use FILL  FILL_490
timestamp 1681620392
transform 1 0 672 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_43
timestamp 1681620392
transform 1 0 680 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_44
timestamp 1681620392
transform 1 0 704 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_45
timestamp 1681620392
transform 1 0 728 0 -1 1770
box -8 -3 32 105
use FILL  FILL_491
timestamp 1681620392
transform 1 0 752 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_46
timestamp 1681620392
transform 1 0 760 0 -1 1770
box -8 -3 32 105
use INVX2  INVX2_149
timestamp 1681620392
transform -1 0 800 0 -1 1770
box -9 -3 26 105
use NAND2X1  NAND2X1_131
timestamp 1681620392
transform 1 0 800 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_132
timestamp 1681620392
transform 1 0 824 0 -1 1770
box -8 -3 32 105
use INVX2  INVX2_150
timestamp 1681620392
transform 1 0 848 0 -1 1770
box -9 -3 26 105
use AOI21X1  AOI21X1_10
timestamp 1681620392
transform -1 0 896 0 -1 1770
box -7 -3 39 105
use NAND2X1  NAND2X1_133
timestamp 1681620392
transform 1 0 896 0 -1 1770
box -8 -3 32 105
use M3_M2  M3_M2_2159
timestamp 1681620392
transform 1 0 932 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_2160
timestamp 1681620392
transform 1 0 996 0 1 1675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_146
timestamp 1681620392
transform 1 0 920 0 -1 1770
box -8 -3 104 105
use M3_M2  M3_M2_2161
timestamp 1681620392
transform 1 0 1052 0 1 1675
box -3 -3 3 3
use OAI22X1  OAI22X1_27
timestamp 1681620392
transform 1 0 1016 0 -1 1770
box -8 -3 46 105
use M3_M2  M3_M2_2162
timestamp 1681620392
transform 1 0 1084 0 1 1675
box -3 -3 3 3
use OAI22X1  OAI22X1_28
timestamp 1681620392
transform -1 0 1096 0 -1 1770
box -8 -3 46 105
use INVX2  INVX2_151
timestamp 1681620392
transform 1 0 1096 0 -1 1770
box -9 -3 26 105
use OAI22X1  OAI22X1_29
timestamp 1681620392
transform -1 0 1152 0 -1 1770
box -8 -3 46 105
use INVX2  INVX2_152
timestamp 1681620392
transform 1 0 1152 0 -1 1770
box -9 -3 26 105
use FILL  FILL_492
timestamp 1681620392
transform 1 0 1168 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_47
timestamp 1681620392
transform 1 0 1176 0 -1 1770
box -8 -3 32 105
use INVX2  INVX2_153
timestamp 1681620392
transform -1 0 1216 0 -1 1770
box -9 -3 26 105
use NOR2X1  NOR2X1_48
timestamp 1681620392
transform -1 0 1240 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_49
timestamp 1681620392
transform 1 0 1240 0 -1 1770
box -8 -3 32 105
use FILL  FILL_493
timestamp 1681620392
transform 1 0 1264 0 -1 1770
box -8 -3 16 105
use AOI21X1  AOI21X1_11
timestamp 1681620392
transform 1 0 1272 0 -1 1770
box -7 -3 39 105
use INVX2  INVX2_154
timestamp 1681620392
transform -1 0 1320 0 -1 1770
box -9 -3 26 105
use NAND2X1  NAND2X1_134
timestamp 1681620392
transform 1 0 1320 0 -1 1770
box -8 -3 32 105
use FILL  FILL_494
timestamp 1681620392
transform 1 0 1344 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_51
timestamp 1681620392
transform 1 0 1352 0 -1 1770
box -8 -3 40 105
use NAND2X1  NAND2X1_135
timestamp 1681620392
transform -1 0 1408 0 -1 1770
box -8 -3 32 105
use FILL  FILL_495
timestamp 1681620392
transform 1 0 1408 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_2163
timestamp 1681620392
transform 1 0 1444 0 1 1675
box -3 -3 3 3
use INVX2  INVX2_155
timestamp 1681620392
transform 1 0 1416 0 -1 1770
box -9 -3 26 105
use FILL  FILL_496
timestamp 1681620392
transform 1 0 1432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_497
timestamp 1681620392
transform 1 0 1440 0 -1 1770
box -8 -3 16 105
use FILL  FILL_498
timestamp 1681620392
transform 1 0 1448 0 -1 1770
box -8 -3 16 105
use FILL  FILL_499
timestamp 1681620392
transform 1 0 1456 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_147
timestamp 1681620392
transform 1 0 1464 0 -1 1770
box -8 -3 104 105
use OAI21X1  OAI21X1_155
timestamp 1681620392
transform -1 0 1592 0 -1 1770
box -8 -3 34 105
use INVX2  INVX2_156
timestamp 1681620392
transform -1 0 1608 0 -1 1770
box -9 -3 26 105
use FILL  FILL_500
timestamp 1681620392
transform 1 0 1608 0 -1 1770
box -8 -3 16 105
use NAND2X1  NAND2X1_136
timestamp 1681620392
transform 1 0 1616 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_137
timestamp 1681620392
transform 1 0 1640 0 -1 1770
box -8 -3 32 105
use FILL  FILL_501
timestamp 1681620392
transform 1 0 1664 0 -1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_156
timestamp 1681620392
transform 1 0 1672 0 -1 1770
box -8 -3 34 105
use FILL  FILL_502
timestamp 1681620392
transform 1 0 1704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_503
timestamp 1681620392
transform 1 0 1712 0 -1 1770
box -8 -3 16 105
use FILL  FILL_504
timestamp 1681620392
transform 1 0 1720 0 -1 1770
box -8 -3 16 105
use FILL  FILL_506
timestamp 1681620392
transform 1 0 1728 0 -1 1770
box -8 -3 16 105
use FILL  FILL_529
timestamp 1681620392
transform 1 0 1736 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_35
timestamp 1681620392
transform -1 0 1784 0 -1 1770
box -8 -3 46 105
use INVX2  INVX2_166
timestamp 1681620392
transform -1 0 1800 0 -1 1770
box -9 -3 26 105
use FILL  FILL_530
timestamp 1681620392
transform 1 0 1800 0 -1 1770
box -8 -3 16 105
use FILL  FILL_531
timestamp 1681620392
transform 1 0 1808 0 -1 1770
box -8 -3 16 105
use FILL  FILL_532
timestamp 1681620392
transform 1 0 1816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_533
timestamp 1681620392
transform 1 0 1824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_534
timestamp 1681620392
transform 1 0 1832 0 -1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_163
timestamp 1681620392
transform -1 0 1872 0 -1 1770
box -8 -3 34 105
use NAND2X1  NAND2X1_142
timestamp 1681620392
transform -1 0 1896 0 -1 1770
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_152
timestamp 1681620392
transform 1 0 1896 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_153
timestamp 1681620392
transform 1 0 1992 0 -1 1770
box -8 -3 104 105
use NAND2X1  NAND2X1_143
timestamp 1681620392
transform 1 0 2088 0 -1 1770
box -8 -3 32 105
use FILL  FILL_535
timestamp 1681620392
transform 1 0 2112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_536
timestamp 1681620392
transform 1 0 2120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_537
timestamp 1681620392
transform 1 0 2128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_538
timestamp 1681620392
transform 1 0 2136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_539
timestamp 1681620392
transform 1 0 2144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_540
timestamp 1681620392
transform 1 0 2152 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_2164
timestamp 1681620392
transform 1 0 2228 0 1 1675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_154
timestamp 1681620392
transform 1 0 2160 0 -1 1770
box -8 -3 104 105
use INVX2  INVX2_167
timestamp 1681620392
transform 1 0 2256 0 -1 1770
box -9 -3 26 105
use FILL  FILL_541
timestamp 1681620392
transform 1 0 2272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_542
timestamp 1681620392
transform 1 0 2280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_543
timestamp 1681620392
transform 1 0 2288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_544
timestamp 1681620392
transform 1 0 2296 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_36
timestamp 1681620392
transform -1 0 2344 0 -1 1770
box -8 -3 46 105
use FILL  FILL_545
timestamp 1681620392
transform 1 0 2344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_546
timestamp 1681620392
transform 1 0 2352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_547
timestamp 1681620392
transform 1 0 2360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_548
timestamp 1681620392
transform 1 0 2368 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_155
timestamp 1681620392
transform 1 0 2376 0 -1 1770
box -8 -3 104 105
use INVX2  INVX2_168
timestamp 1681620392
transform -1 0 2488 0 -1 1770
box -9 -3 26 105
use FILL  FILL_549
timestamp 1681620392
transform 1 0 2488 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_156
timestamp 1681620392
transform 1 0 2496 0 -1 1770
box -8 -3 104 105
use OAI21X1  OAI21X1_164
timestamp 1681620392
transform -1 0 2624 0 -1 1770
box -8 -3 34 105
use INVX2  INVX2_169
timestamp 1681620392
transform 1 0 2624 0 -1 1770
box -9 -3 26 105
use FILL  FILL_550
timestamp 1681620392
transform 1 0 2640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_551
timestamp 1681620392
transform 1 0 2648 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_157
timestamp 1681620392
transform -1 0 2752 0 -1 1770
box -8 -3 104 105
use FILL  FILL_552
timestamp 1681620392
transform 1 0 2752 0 -1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_165
timestamp 1681620392
transform 1 0 2760 0 -1 1770
box -8 -3 34 105
use INVX2  INVX2_170
timestamp 1681620392
transform 1 0 2792 0 -1 1770
box -9 -3 26 105
use FILL  FILL_553
timestamp 1681620392
transform 1 0 2808 0 -1 1770
box -8 -3 16 105
use FILL  FILL_554
timestamp 1681620392
transform 1 0 2816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_555
timestamp 1681620392
transform 1 0 2824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_556
timestamp 1681620392
transform 1 0 2832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_557
timestamp 1681620392
transform 1 0 2840 0 -1 1770
box -8 -3 16 105
use NAND2X1  NAND2X1_144
timestamp 1681620392
transform 1 0 2848 0 -1 1770
box -8 -3 32 105
use OAI21X1  OAI21X1_166
timestamp 1681620392
transform 1 0 2872 0 -1 1770
box -8 -3 34 105
use INVX2  INVX2_171
timestamp 1681620392
transform 1 0 2904 0 -1 1770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_158
timestamp 1681620392
transform 1 0 2920 0 -1 1770
box -8 -3 104 105
use Project_Top_VIA0  Project_Top_VIA0_27
timestamp 1681620392
transform 1 0 3067 0 1 1670
box -10 -3 10 3
use M2_M1  M2_M1_2580
timestamp 1681620392
transform 1 0 132 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2257
timestamp 1681620392
transform 1 0 148 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2219
timestamp 1681620392
transform 1 0 180 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2220
timestamp 1681620392
transform 1 0 204 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2581
timestamp 1681620392
transform 1 0 164 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2582
timestamp 1681620392
transform 1 0 180 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2258
timestamp 1681620392
transform 1 0 188 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_2583
timestamp 1681620392
transform 1 0 196 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2664
timestamp 1681620392
transform 1 0 84 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2276
timestamp 1681620392
transform 1 0 164 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_2665
timestamp 1681620392
transform 1 0 172 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2277
timestamp 1681620392
transform 1 0 180 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_2666
timestamp 1681620392
transform 1 0 188 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2298
timestamp 1681620392
transform 1 0 84 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2299
timestamp 1681620392
transform 1 0 108 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2300
timestamp 1681620392
transform 1 0 132 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2323
timestamp 1681620392
transform 1 0 84 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2324
timestamp 1681620392
transform 1 0 124 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2301
timestamp 1681620392
transform 1 0 188 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_2667
timestamp 1681620392
transform 1 0 212 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2668
timestamp 1681620392
transform 1 0 220 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2302
timestamp 1681620392
transform 1 0 212 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2173
timestamp 1681620392
transform 1 0 244 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2221
timestamp 1681620392
transform 1 0 236 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2584
timestamp 1681620392
transform 1 0 228 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2278
timestamp 1681620392
transform 1 0 228 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_2669
timestamp 1681620392
transform 1 0 236 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2174
timestamp 1681620392
transform 1 0 284 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2190
timestamp 1681620392
transform 1 0 260 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_2670
timestamp 1681620392
transform 1 0 252 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2303
timestamp 1681620392
transform 1 0 252 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2222
timestamp 1681620392
transform 1 0 284 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2585
timestamp 1681620392
transform 1 0 268 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2586
timestamp 1681620392
transform 1 0 284 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2279
timestamp 1681620392
transform 1 0 268 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2223
timestamp 1681620392
transform 1 0 324 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2587
timestamp 1681620392
transform 1 0 308 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2588
timestamp 1681620392
transform 1 0 324 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2671
timestamp 1681620392
transform 1 0 276 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2672
timestamp 1681620392
transform 1 0 292 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2673
timestamp 1681620392
transform 1 0 300 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2674
timestamp 1681620392
transform 1 0 316 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2280
timestamp 1681620392
transform 1 0 324 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2191
timestamp 1681620392
transform 1 0 388 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_2589
timestamp 1681620392
transform 1 0 388 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2675
timestamp 1681620392
transform 1 0 332 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2676
timestamp 1681620392
transform 1 0 348 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2677
timestamp 1681620392
transform 1 0 436 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2304
timestamp 1681620392
transform 1 0 300 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2305
timestamp 1681620392
transform 1 0 316 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2306
timestamp 1681620392
transform 1 0 388 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2307
timestamp 1681620392
transform 1 0 436 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2165
timestamp 1681620392
transform 1 0 556 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2175
timestamp 1681620392
transform 1 0 572 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2224
timestamp 1681620392
transform 1 0 540 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2590
timestamp 1681620392
transform 1 0 500 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2591
timestamp 1681620392
transform 1 0 540 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2592
timestamp 1681620392
transform 1 0 556 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2593
timestamp 1681620392
transform 1 0 572 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2678
timestamp 1681620392
transform 1 0 460 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2679
timestamp 1681620392
transform 1 0 548 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2308
timestamp 1681620392
transform 1 0 460 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2281
timestamp 1681620392
transform 1 0 556 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_2680
timestamp 1681620392
transform 1 0 564 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2681
timestamp 1681620392
transform 1 0 580 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2682
timestamp 1681620392
transform 1 0 588 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2309
timestamp 1681620392
transform 1 0 580 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2225
timestamp 1681620392
transform 1 0 604 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2594
timestamp 1681620392
transform 1 0 604 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2282
timestamp 1681620392
transform 1 0 628 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_2683
timestamp 1681620392
transform 1 0 636 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2750
timestamp 1681620392
transform 1 0 628 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_2310
timestamp 1681620392
transform 1 0 636 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_2595
timestamp 1681620392
transform 1 0 652 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2596
timestamp 1681620392
transform 1 0 668 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2192
timestamp 1681620392
transform 1 0 684 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_2552
timestamp 1681620392
transform 1 0 684 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2684
timestamp 1681620392
transform 1 0 676 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2685
timestamp 1681620392
transform 1 0 700 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2325
timestamp 1681620392
transform 1 0 700 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2167
timestamp 1681620392
transform 1 0 716 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_2597
timestamp 1681620392
transform 1 0 716 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2259
timestamp 1681620392
transform 1 0 732 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2283
timestamp 1681620392
transform 1 0 716 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2260
timestamp 1681620392
transform 1 0 756 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_2686
timestamp 1681620392
transform 1 0 724 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2687
timestamp 1681620392
transform 1 0 732 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2326
timestamp 1681620392
transform 1 0 724 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2284
timestamp 1681620392
transform 1 0 748 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_2688
timestamp 1681620392
transform 1 0 756 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2751
timestamp 1681620392
transform 1 0 748 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_2598
timestamp 1681620392
transform 1 0 780 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2193
timestamp 1681620392
transform 1 0 796 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_2553
timestamp 1681620392
transform 1 0 796 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2689
timestamp 1681620392
transform 1 0 804 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2311
timestamp 1681620392
transform 1 0 804 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2226
timestamp 1681620392
transform 1 0 828 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2545
timestamp 1681620392
transform 1 0 860 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2554
timestamp 1681620392
transform 1 0 844 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2555
timestamp 1681620392
transform 1 0 852 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2599
timestamp 1681620392
transform 1 0 828 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2600
timestamp 1681620392
transform 1 0 836 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2690
timestamp 1681620392
transform 1 0 820 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2227
timestamp 1681620392
transform 1 0 868 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2556
timestamp 1681620392
transform 1 0 876 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2557
timestamp 1681620392
transform 1 0 884 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2601
timestamp 1681620392
transform 1 0 868 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2327
timestamp 1681620392
transform 1 0 884 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2176
timestamp 1681620392
transform 1 0 908 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2194
timestamp 1681620392
transform 1 0 900 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_2546
timestamp 1681620392
transform 1 0 924 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2558
timestamp 1681620392
transform 1 0 908 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_2228
timestamp 1681620392
transform 1 0 916 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2195
timestamp 1681620392
transform 1 0 940 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_2559
timestamp 1681620392
transform 1 0 932 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2560
timestamp 1681620392
transform 1 0 940 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2602
timestamp 1681620392
transform 1 0 900 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2603
timestamp 1681620392
transform 1 0 916 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2691
timestamp 1681620392
transform 1 0 900 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2177
timestamp 1681620392
transform 1 0 956 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_2547
timestamp 1681620392
transform 1 0 964 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2561
timestamp 1681620392
transform 1 0 972 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2604
timestamp 1681620392
transform 1 0 956 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2178
timestamp 1681620392
transform 1 0 1012 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2179
timestamp 1681620392
transform 1 0 1044 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2166
timestamp 1681620392
transform 1 0 1092 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2196
timestamp 1681620392
transform 1 0 1108 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2229
timestamp 1681620392
transform 1 0 1076 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2605
timestamp 1681620392
transform 1 0 1036 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2606
timestamp 1681620392
transform 1 0 1076 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2607
timestamp 1681620392
transform 1 0 1092 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2608
timestamp 1681620392
transform 1 0 1108 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2168
timestamp 1681620392
transform 1 0 1148 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2197
timestamp 1681620392
transform 1 0 1140 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2230
timestamp 1681620392
transform 1 0 1140 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2609
timestamp 1681620392
transform 1 0 1132 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2610
timestamp 1681620392
transform 1 0 1140 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2692
timestamp 1681620392
transform 1 0 996 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2693
timestamp 1681620392
transform 1 0 1084 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2694
timestamp 1681620392
transform 1 0 1100 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2695
timestamp 1681620392
transform 1 0 1124 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2285
timestamp 1681620392
transform 1 0 1132 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2286
timestamp 1681620392
transform 1 0 1156 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_2696
timestamp 1681620392
transform 1 0 1164 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2752
timestamp 1681620392
transform 1 0 1156 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_2328
timestamp 1681620392
transform 1 0 1164 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2180
timestamp 1681620392
transform 1 0 1180 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_2611
timestamp 1681620392
transform 1 0 1180 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2697
timestamp 1681620392
transform 1 0 1188 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2753
timestamp 1681620392
transform 1 0 1196 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_2612
timestamp 1681620392
transform 1 0 1212 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2613
timestamp 1681620392
transform 1 0 1244 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2698
timestamp 1681620392
transform 1 0 1236 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2198
timestamp 1681620392
transform 1 0 1268 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2261
timestamp 1681620392
transform 1 0 1260 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_2699
timestamp 1681620392
transform 1 0 1252 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2700
timestamp 1681620392
transform 1 0 1260 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2329
timestamp 1681620392
transform 1 0 1252 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2330
timestamp 1681620392
transform 1 0 1268 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2181
timestamp 1681620392
transform 1 0 1324 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_2548
timestamp 1681620392
transform 1 0 1316 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2562
timestamp 1681620392
transform 1 0 1292 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_2231
timestamp 1681620392
transform 1 0 1300 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2199
timestamp 1681620392
transform 1 0 1332 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_2563
timestamp 1681620392
transform 1 0 1308 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2564
timestamp 1681620392
transform 1 0 1324 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2565
timestamp 1681620392
transform 1 0 1332 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2614
timestamp 1681620392
transform 1 0 1284 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2615
timestamp 1681620392
transform 1 0 1308 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2616
timestamp 1681620392
transform 1 0 1332 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2701
timestamp 1681620392
transform 1 0 1292 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2331
timestamp 1681620392
transform 1 0 1332 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2262
timestamp 1681620392
transform 1 0 1348 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_2702
timestamp 1681620392
transform 1 0 1348 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2182
timestamp 1681620392
transform 1 0 1364 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2200
timestamp 1681620392
transform 1 0 1388 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2232
timestamp 1681620392
transform 1 0 1380 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2566
timestamp 1681620392
transform 1 0 1388 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_2201
timestamp 1681620392
transform 1 0 1420 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_2617
timestamp 1681620392
transform 1 0 1380 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2703
timestamp 1681620392
transform 1 0 1372 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2263
timestamp 1681620392
transform 1 0 1388 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_2618
timestamp 1681620392
transform 1 0 1396 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2264
timestamp 1681620392
transform 1 0 1404 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_2619
timestamp 1681620392
transform 1 0 1420 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2620
timestamp 1681620392
transform 1 0 1428 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2704
timestamp 1681620392
transform 1 0 1388 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2287
timestamp 1681620392
transform 1 0 1420 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_2754
timestamp 1681620392
transform 1 0 1420 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_2233
timestamp 1681620392
transform 1 0 1436 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2621
timestamp 1681620392
transform 1 0 1444 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2705
timestamp 1681620392
transform 1 0 1436 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2288
timestamp 1681620392
transform 1 0 1444 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2234
timestamp 1681620392
transform 1 0 1460 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2265
timestamp 1681620392
transform 1 0 1468 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_2706
timestamp 1681620392
transform 1 0 1468 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2567
timestamp 1681620392
transform 1 0 1508 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_2183
timestamp 1681620392
transform 1 0 1572 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2202
timestamp 1681620392
transform 1 0 1548 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2203
timestamp 1681620392
transform 1 0 1564 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_2549
timestamp 1681620392
transform 1 0 1572 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_2204
timestamp 1681620392
transform 1 0 1596 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2235
timestamp 1681620392
transform 1 0 1540 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2236
timestamp 1681620392
transform 1 0 1556 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2568
timestamp 1681620392
transform 1 0 1564 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_2237
timestamp 1681620392
transform 1 0 1572 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2569
timestamp 1681620392
transform 1 0 1588 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2622
timestamp 1681620392
transform 1 0 1532 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2707
timestamp 1681620392
transform 1 0 1516 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2332
timestamp 1681620392
transform 1 0 1516 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_2623
timestamp 1681620392
transform 1 0 1556 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2624
timestamp 1681620392
transform 1 0 1572 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2708
timestamp 1681620392
transform 1 0 1540 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2333
timestamp 1681620392
transform 1 0 1540 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2266
timestamp 1681620392
transform 1 0 1580 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_2625
timestamp 1681620392
transform 1 0 1596 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2267
timestamp 1681620392
transform 1 0 1604 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2184
timestamp 1681620392
transform 1 0 1652 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_2550
timestamp 1681620392
transform 1 0 1652 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_2238
timestamp 1681620392
transform 1 0 1636 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2570
timestamp 1681620392
transform 1 0 1652 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2626
timestamp 1681620392
transform 1 0 1628 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2709
timestamp 1681620392
transform 1 0 1604 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2289
timestamp 1681620392
transform 1 0 1628 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2239
timestamp 1681620392
transform 1 0 1660 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2571
timestamp 1681620392
transform 1 0 1684 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2627
timestamp 1681620392
transform 1 0 1644 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2628
timestamp 1681620392
transform 1 0 1660 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2710
timestamp 1681620392
transform 1 0 1636 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2312
timestamp 1681620392
transform 1 0 1612 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_2755
timestamp 1681620392
transform 1 0 1620 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_2756
timestamp 1681620392
transform 1 0 1628 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_2313
timestamp 1681620392
transform 1 0 1636 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2334
timestamp 1681620392
transform 1 0 1620 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2205
timestamp 1681620392
transform 1 0 1700 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2169
timestamp 1681620392
transform 1 0 1820 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2170
timestamp 1681620392
transform 1 0 1940 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2240
timestamp 1681620392
transform 1 0 1916 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2629
timestamp 1681620392
transform 1 0 1700 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2630
timestamp 1681620392
transform 1 0 1764 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2631
timestamp 1681620392
transform 1 0 1796 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2632
timestamp 1681620392
transform 1 0 1836 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2633
timestamp 1681620392
transform 1 0 1892 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2634
timestamp 1681620392
transform 1 0 1900 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2711
timestamp 1681620392
transform 1 0 1700 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2712
timestamp 1681620392
transform 1 0 1716 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2290
timestamp 1681620392
transform 1 0 1740 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2314
timestamp 1681620392
transform 1 0 1716 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2315
timestamp 1681620392
transform 1 0 1788 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_2713
timestamp 1681620392
transform 1 0 1812 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2316
timestamp 1681620392
transform 1 0 1812 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2317
timestamp 1681620392
transform 1 0 1852 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_2635
timestamp 1681620392
transform 1 0 1924 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2241
timestamp 1681620392
transform 1 0 1964 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2206
timestamp 1681620392
transform 1 0 2020 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2242
timestamp 1681620392
transform 1 0 1996 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2636
timestamp 1681620392
transform 1 0 1964 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2714
timestamp 1681620392
transform 1 0 1916 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2715
timestamp 1681620392
transform 1 0 1940 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2716
timestamp 1681620392
transform 1 0 1948 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2318
timestamp 1681620392
transform 1 0 1948 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2268
timestamp 1681620392
transform 1 0 1988 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_2637
timestamp 1681620392
transform 1 0 1996 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2717
timestamp 1681620392
transform 1 0 1988 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2243
timestamp 1681620392
transform 1 0 2028 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2244
timestamp 1681620392
transform 1 0 2060 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2638
timestamp 1681620392
transform 1 0 2028 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2639
timestamp 1681620392
transform 1 0 2044 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2640
timestamp 1681620392
transform 1 0 2060 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2718
timestamp 1681620392
transform 1 0 2012 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2719
timestamp 1681620392
transform 1 0 2020 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2720
timestamp 1681620392
transform 1 0 2036 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2291
timestamp 1681620392
transform 1 0 2044 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_2721
timestamp 1681620392
transform 1 0 2052 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2722
timestamp 1681620392
transform 1 0 2076 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2207
timestamp 1681620392
transform 1 0 2108 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_2723
timestamp 1681620392
transform 1 0 2100 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2208
timestamp 1681620392
transform 1 0 2148 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_2641
timestamp 1681620392
transform 1 0 2124 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2292
timestamp 1681620392
transform 1 0 2124 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_2724
timestamp 1681620392
transform 1 0 2132 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2725
timestamp 1681620392
transform 1 0 2148 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2642
timestamp 1681620392
transform 1 0 2164 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2209
timestamp 1681620392
transform 1 0 2204 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_2643
timestamp 1681620392
transform 1 0 2180 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2726
timestamp 1681620392
transform 1 0 2172 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2335
timestamp 1681620392
transform 1 0 2164 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2293
timestamp 1681620392
transform 1 0 2180 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2245
timestamp 1681620392
transform 1 0 2212 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2644
timestamp 1681620392
transform 1 0 2212 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2727
timestamp 1681620392
transform 1 0 2188 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2728
timestamp 1681620392
transform 1 0 2204 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2336
timestamp 1681620392
transform 1 0 2188 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2210
timestamp 1681620392
transform 1 0 2340 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2246
timestamp 1681620392
transform 1 0 2276 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2247
timestamp 1681620392
transform 1 0 2300 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2248
timestamp 1681620392
transform 1 0 2324 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2269
timestamp 1681620392
transform 1 0 2252 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_2645
timestamp 1681620392
transform 1 0 2300 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2729
timestamp 1681620392
transform 1 0 2252 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2294
timestamp 1681620392
transform 1 0 2316 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2211
timestamp 1681620392
transform 1 0 2380 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2249
timestamp 1681620392
transform 1 0 2372 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2250
timestamp 1681620392
transform 1 0 2428 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2646
timestamp 1681620392
transform 1 0 2348 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2647
timestamp 1681620392
transform 1 0 2364 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2648
timestamp 1681620392
transform 1 0 2380 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2270
timestamp 1681620392
transform 1 0 2388 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_2649
timestamp 1681620392
transform 1 0 2428 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2271
timestamp 1681620392
transform 1 0 2476 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_2650
timestamp 1681620392
transform 1 0 2484 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2730
timestamp 1681620392
transform 1 0 2356 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2295
timestamp 1681620392
transform 1 0 2364 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_2731
timestamp 1681620392
transform 1 0 2372 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2732
timestamp 1681620392
transform 1 0 2388 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2733
timestamp 1681620392
transform 1 0 2404 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2337
timestamp 1681620392
transform 1 0 2372 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_2651
timestamp 1681620392
transform 1 0 2516 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2734
timestamp 1681620392
transform 1 0 2500 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2735
timestamp 1681620392
transform 1 0 2508 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2757
timestamp 1681620392
transform 1 0 2492 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_2338
timestamp 1681620392
transform 1 0 2436 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2296
timestamp 1681620392
transform 1 0 2516 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2339
timestamp 1681620392
transform 1 0 2508 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_2652
timestamp 1681620392
transform 1 0 2548 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2736
timestamp 1681620392
transform 1 0 2564 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2251
timestamp 1681620392
transform 1 0 2588 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2212
timestamp 1681620392
transform 1 0 2628 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_2572
timestamp 1681620392
transform 1 0 2612 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2573
timestamp 1681620392
transform 1 0 2628 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2653
timestamp 1681620392
transform 1 0 2588 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2654
timestamp 1681620392
transform 1 0 2604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2737
timestamp 1681620392
transform 1 0 2580 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2252
timestamp 1681620392
transform 1 0 2636 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2655
timestamp 1681620392
transform 1 0 2636 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2297
timestamp 1681620392
transform 1 0 2644 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2185
timestamp 1681620392
transform 1 0 2668 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_2574
timestamp 1681620392
transform 1 0 2684 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2656
timestamp 1681620392
transform 1 0 2668 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2738
timestamp 1681620392
transform 1 0 2660 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2213
timestamp 1681620392
transform 1 0 2700 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_2657
timestamp 1681620392
transform 1 0 2700 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_2171
timestamp 1681620392
transform 1 0 2756 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2214
timestamp 1681620392
transform 1 0 2748 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2186
timestamp 1681620392
transform 1 0 2772 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2215
timestamp 1681620392
transform 1 0 2764 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_2575
timestamp 1681620392
transform 1 0 2756 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_2272
timestamp 1681620392
transform 1 0 2724 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2273
timestamp 1681620392
transform 1 0 2740 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_2739
timestamp 1681620392
transform 1 0 2700 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2740
timestamp 1681620392
transform 1 0 2708 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2319
timestamp 1681620392
transform 1 0 2700 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_2741
timestamp 1681620392
transform 1 0 2732 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2742
timestamp 1681620392
transform 1 0 2740 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2320
timestamp 1681620392
transform 1 0 2740 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2187
timestamp 1681620392
transform 1 0 2804 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2216
timestamp 1681620392
transform 1 0 2788 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_2576
timestamp 1681620392
transform 1 0 2788 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_2253
timestamp 1681620392
transform 1 0 2796 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2188
timestamp 1681620392
transform 1 0 2844 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_2551
timestamp 1681620392
transform 1 0 2844 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_2217
timestamp 1681620392
transform 1 0 2852 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_2577
timestamp 1681620392
transform 1 0 2820 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_2274
timestamp 1681620392
transform 1 0 2788 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_2658
timestamp 1681620392
transform 1 0 2804 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2743
timestamp 1681620392
transform 1 0 2788 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2321
timestamp 1681620392
transform 1 0 2788 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2254
timestamp 1681620392
transform 1 0 2828 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2578
timestamp 1681620392
transform 1 0 2852 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_2275
timestamp 1681620392
transform 1 0 2828 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2172
timestamp 1681620392
transform 1 0 2868 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2218
timestamp 1681620392
transform 1 0 2876 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_2579
timestamp 1681620392
transform 1 0 2868 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2659
timestamp 1681620392
transform 1 0 2860 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2744
timestamp 1681620392
transform 1 0 2812 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2745
timestamp 1681620392
transform 1 0 2836 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2746
timestamp 1681620392
transform 1 0 2852 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2322
timestamp 1681620392
transform 1 0 2852 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_2660
timestamp 1681620392
transform 1 0 2876 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2661
timestamp 1681620392
transform 1 0 2892 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2747
timestamp 1681620392
transform 1 0 2892 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2189
timestamp 1681620392
transform 1 0 2980 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2255
timestamp 1681620392
transform 1 0 2916 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2256
timestamp 1681620392
transform 1 0 3012 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_2662
timestamp 1681620392
transform 1 0 2956 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2663
timestamp 1681620392
transform 1 0 3012 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2748
timestamp 1681620392
transform 1 0 2916 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2749
timestamp 1681620392
transform 1 0 2932 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_2340
timestamp 1681620392
transform 1 0 2932 0 1 1585
box -3 -3 3 3
use Project_Top_VIA0  Project_Top_VIA0_28
timestamp 1681620392
transform 1 0 48 0 1 1570
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_159
timestamp 1681620392
transform 1 0 72 0 1 1570
box -8 -3 104 105
use OAI22X1  OAI22X1_37
timestamp 1681620392
transform 1 0 168 0 1 1570
box -8 -3 46 105
use FILL  FILL_558
timestamp 1681620392
transform 1 0 208 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_172
timestamp 1681620392
transform 1 0 216 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_173
timestamp 1681620392
transform 1 0 232 0 1 1570
box -9 -3 26 105
use FILL  FILL_559
timestamp 1681620392
transform 1 0 248 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_38
timestamp 1681620392
transform -1 0 296 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_39
timestamp 1681620392
transform -1 0 336 0 1 1570
box -8 -3 46 105
use INVX2  INVX2_174
timestamp 1681620392
transform -1 0 352 0 1 1570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_160
timestamp 1681620392
transform -1 0 448 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_161
timestamp 1681620392
transform 1 0 448 0 1 1570
box -8 -3 104 105
use OAI22X1  OAI22X1_40
timestamp 1681620392
transform -1 0 584 0 1 1570
box -8 -3 46 105
use INVX2  INVX2_175
timestamp 1681620392
transform 1 0 584 0 1 1570
box -9 -3 26 105
use FILL  FILL_560
timestamp 1681620392
transform 1 0 600 0 1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_50
timestamp 1681620392
transform -1 0 632 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_51
timestamp 1681620392
transform 1 0 632 0 1 1570
box -8 -3 32 105
use FILL  FILL_561
timestamp 1681620392
transform 1 0 656 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_2341
timestamp 1681620392
transform 1 0 676 0 1 1575
box -3 -3 3 3
use FILL  FILL_580
timestamp 1681620392
transform 1 0 664 0 1 1570
box -8 -3 16 105
use FILL  FILL_582
timestamp 1681620392
transform 1 0 672 0 1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_146
timestamp 1681620392
transform -1 0 704 0 1 1570
box -8 -3 32 105
use INVX2  INVX2_179
timestamp 1681620392
transform 1 0 704 0 1 1570
box -9 -3 26 105
use AOI21X1  AOI21X1_13
timestamp 1681620392
transform 1 0 720 0 1 1570
box -7 -3 39 105
use FILL  FILL_583
timestamp 1681620392
transform 1 0 752 0 1 1570
box -8 -3 16 105
use FILL  FILL_588
timestamp 1681620392
transform 1 0 760 0 1 1570
box -8 -3 16 105
use FILL  FILL_590
timestamp 1681620392
transform 1 0 768 0 1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_148
timestamp 1681620392
transform 1 0 776 0 1 1570
box -8 -3 32 105
use FILL  FILL_591
timestamp 1681620392
transform 1 0 800 0 1 1570
box -8 -3 16 105
use FILL  FILL_594
timestamp 1681620392
transform 1 0 808 0 1 1570
box -8 -3 16 105
use FILL  FILL_596
timestamp 1681620392
transform 1 0 816 0 1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_150
timestamp 1681620392
transform 1 0 824 0 1 1570
box -8 -3 32 105
use NAND3X1  NAND3X1_53
timestamp 1681620392
transform -1 0 880 0 1 1570
box -8 -3 40 105
use M3_M2  M3_M2_2342
timestamp 1681620392
transform 1 0 900 0 1 1575
box -3 -3 3 3
use NAND2X1  NAND2X1_151
timestamp 1681620392
transform -1 0 904 0 1 1570
box -8 -3 32 105
use NAND3X1  NAND3X1_54
timestamp 1681620392
transform 1 0 904 0 1 1570
box -8 -3 40 105
use FILL  FILL_598
timestamp 1681620392
transform 1 0 936 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_55
timestamp 1681620392
transform 1 0 944 0 1 1570
box -8 -3 40 105
use FILL  FILL_599
timestamp 1681620392
transform 1 0 976 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_164
timestamp 1681620392
transform 1 0 984 0 1 1570
box -8 -3 104 105
use OAI22X1  OAI22X1_42
timestamp 1681620392
transform -1 0 1120 0 1 1570
box -8 -3 46 105
use INVX2  INVX2_180
timestamp 1681620392
transform 1 0 1120 0 1 1570
box -9 -3 26 105
use NOR2X1  NOR2X1_58
timestamp 1681620392
transform -1 0 1160 0 1 1570
box -8 -3 32 105
use M3_M2  M3_M2_2343
timestamp 1681620392
transform 1 0 1188 0 1 1575
box -3 -3 3 3
use NOR2X1  NOR2X1_59
timestamp 1681620392
transform 1 0 1160 0 1 1570
box -8 -3 32 105
use FILL  FILL_600
timestamp 1681620392
transform 1 0 1184 0 1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_62
timestamp 1681620392
transform 1 0 1192 0 1 1570
box -8 -3 32 105
use FILL  FILL_619
timestamp 1681620392
transform 1 0 1216 0 1 1570
box -8 -3 16 105
use FILL  FILL_620
timestamp 1681620392
transform 1 0 1224 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_2344
timestamp 1681620392
transform 1 0 1260 0 1 1575
box -3 -3 3 3
use NAND2X1  NAND2X1_155
timestamp 1681620392
transform -1 0 1256 0 1 1570
box -8 -3 32 105
use FILL  FILL_621
timestamp 1681620392
transform 1 0 1256 0 1 1570
box -8 -3 16 105
use FILL  FILL_622
timestamp 1681620392
transform 1 0 1264 0 1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_158
timestamp 1681620392
transform 1 0 1272 0 1 1570
box -8 -3 32 105
use NAND3X1  NAND3X1_57
timestamp 1681620392
transform 1 0 1296 0 1 1570
box -8 -3 40 105
use NAND2X1  NAND2X1_159
timestamp 1681620392
transform -1 0 1352 0 1 1570
box -8 -3 32 105
use FILL  FILL_624
timestamp 1681620392
transform 1 0 1352 0 1 1570
box -8 -3 16 105
use FILL  FILL_625
timestamp 1681620392
transform 1 0 1360 0 1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_160
timestamp 1681620392
transform 1 0 1368 0 1 1570
box -8 -3 32 105
use AOI21X1  AOI21X1_15
timestamp 1681620392
transform 1 0 1392 0 1 1570
box -7 -3 39 105
use INVX2  INVX2_183
timestamp 1681620392
transform -1 0 1440 0 1 1570
box -9 -3 26 105
use FILL  FILL_626
timestamp 1681620392
transform 1 0 1440 0 1 1570
box -8 -3 16 105
use FILL  FILL_635
timestamp 1681620392
transform 1 0 1448 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_184
timestamp 1681620392
transform -1 0 1472 0 1 1570
box -9 -3 26 105
use FILL  FILL_636
timestamp 1681620392
transform 1 0 1472 0 1 1570
box -8 -3 16 105
use FILL  FILL_637
timestamp 1681620392
transform 1 0 1480 0 1 1570
box -8 -3 16 105
use FILL  FILL_639
timestamp 1681620392
transform 1 0 1488 0 1 1570
box -8 -3 16 105
use FILL  FILL_641
timestamp 1681620392
transform 1 0 1496 0 1 1570
box -8 -3 16 105
use FILL  FILL_643
timestamp 1681620392
transform 1 0 1504 0 1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_168
timestamp 1681620392
transform -1 0 1544 0 1 1570
box -8 -3 34 105
use INVX2  INVX2_185
timestamp 1681620392
transform 1 0 1544 0 1 1570
box -9 -3 26 105
use NAND3X1  NAND3X1_60
timestamp 1681620392
transform 1 0 1560 0 1 1570
box -8 -3 40 105
use M3_M2  M3_M2_2345
timestamp 1681620392
transform 1 0 1620 0 1 1575
box -3 -3 3 3
use AOI21X1  AOI21X1_17
timestamp 1681620392
transform 1 0 1592 0 1 1570
box -7 -3 39 105
use M3_M2  M3_M2_2346
timestamp 1681620392
transform 1 0 1652 0 1 1575
box -3 -3 3 3
use NOR2X1  NOR2X1_63
timestamp 1681620392
transform 1 0 1624 0 1 1570
box -8 -3 32 105
use NAND3X1  NAND3X1_61
timestamp 1681620392
transform 1 0 1648 0 1 1570
box -8 -3 40 105
use NAND2X1  NAND2X1_163
timestamp 1681620392
transform -1 0 1704 0 1 1570
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_165
timestamp 1681620392
transform 1 0 1704 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_166
timestamp 1681620392
transform 1 0 1800 0 1 1570
box -8 -3 104 105
use BUFX2  BUFX2_18
timestamp 1681620392
transform 1 0 1896 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_19
timestamp 1681620392
transform 1 0 1920 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_20
timestamp 1681620392
transform -1 0 1968 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_21
timestamp 1681620392
transform 1 0 1968 0 1 1570
box -5 -3 28 105
use M3_M2  M3_M2_2347
timestamp 1681620392
transform 1 0 2044 0 1 1575
box -3 -3 3 3
use BUFX2  BUFX2_22
timestamp 1681620392
transform 1 0 1992 0 1 1570
box -5 -3 28 105
use OAI22X1  OAI22X1_43
timestamp 1681620392
transform 1 0 2016 0 1 1570
box -8 -3 46 105
use INVX2  INVX2_186
timestamp 1681620392
transform -1 0 2072 0 1 1570
box -9 -3 26 105
use FILL  FILL_644
timestamp 1681620392
transform 1 0 2072 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_2348
timestamp 1681620392
transform 1 0 2100 0 1 1575
box -3 -3 3 3
use FILL  FILL_645
timestamp 1681620392
transform 1 0 2080 0 1 1570
box -8 -3 16 105
use FILL  FILL_646
timestamp 1681620392
transform 1 0 2088 0 1 1570
box -8 -3 16 105
use FILL  FILL_647
timestamp 1681620392
transform 1 0 2096 0 1 1570
box -8 -3 16 105
use FILL  FILL_648
timestamp 1681620392
transform 1 0 2104 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_44
timestamp 1681620392
transform -1 0 2152 0 1 1570
box -8 -3 46 105
use FILL  FILL_649
timestamp 1681620392
transform 1 0 2152 0 1 1570
box -8 -3 16 105
use FILL  FILL_650
timestamp 1681620392
transform 1 0 2160 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_45
timestamp 1681620392
transform -1 0 2208 0 1 1570
box -8 -3 46 105
use FILL  FILL_651
timestamp 1681620392
transform 1 0 2208 0 1 1570
box -8 -3 16 105
use FILL  FILL_652
timestamp 1681620392
transform 1 0 2216 0 1 1570
box -8 -3 16 105
use FILL  FILL_653
timestamp 1681620392
transform 1 0 2224 0 1 1570
box -8 -3 16 105
use FILL  FILL_654
timestamp 1681620392
transform 1 0 2232 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_2349
timestamp 1681620392
transform 1 0 2252 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_167
timestamp 1681620392
transform 1 0 2240 0 1 1570
box -8 -3 104 105
use INVX2  INVX2_187
timestamp 1681620392
transform 1 0 2336 0 1 1570
box -9 -3 26 105
use OAI22X1  OAI22X1_46
timestamp 1681620392
transform -1 0 2392 0 1 1570
box -8 -3 46 105
use M3_M2  M3_M2_2350
timestamp 1681620392
transform 1 0 2404 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_168
timestamp 1681620392
transform 1 0 2392 0 1 1570
box -8 -3 104 105
use NOR2X1  NOR2X1_64
timestamp 1681620392
transform 1 0 2488 0 1 1570
box -8 -3 32 105
use FILL  FILL_655
timestamp 1681620392
transform 1 0 2512 0 1 1570
box -8 -3 16 105
use BUFX2  BUFX2_23
timestamp 1681620392
transform -1 0 2544 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_24
timestamp 1681620392
transform 1 0 2544 0 1 1570
box -5 -3 28 105
use FILL  FILL_656
timestamp 1681620392
transform 1 0 2568 0 1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_169
timestamp 1681620392
transform 1 0 2576 0 1 1570
box -8 -3 34 105
use NAND2X1  NAND2X1_164
timestamp 1681620392
transform 1 0 2608 0 1 1570
box -8 -3 32 105
use FILL  FILL_657
timestamp 1681620392
transform 1 0 2632 0 1 1570
box -8 -3 16 105
use FILL  FILL_658
timestamp 1681620392
transform 1 0 2640 0 1 1570
box -8 -3 16 105
use FILL  FILL_659
timestamp 1681620392
transform 1 0 2648 0 1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_170
timestamp 1681620392
transform 1 0 2656 0 1 1570
box -8 -3 34 105
use FILL  FILL_660
timestamp 1681620392
transform 1 0 2688 0 1 1570
box -8 -3 16 105
use FILL  FILL_661
timestamp 1681620392
transform 1 0 2696 0 1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_171
timestamp 1681620392
transform 1 0 2704 0 1 1570
box -8 -3 34 105
use NAND2X1  NAND2X1_165
timestamp 1681620392
transform 1 0 2736 0 1 1570
box -8 -3 32 105
use FILL  FILL_662
timestamp 1681620392
transform 1 0 2760 0 1 1570
box -8 -3 16 105
use FILL  FILL_663
timestamp 1681620392
transform 1 0 2768 0 1 1570
box -8 -3 16 105
use FILL  FILL_664
timestamp 1681620392
transform 1 0 2776 0 1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_172
timestamp 1681620392
transform -1 0 2816 0 1 1570
box -8 -3 34 105
use NAND3X1  NAND3X1_62
timestamp 1681620392
transform -1 0 2848 0 1 1570
box -8 -3 40 105
use NAND2X1  NAND2X1_166
timestamp 1681620392
transform 1 0 2848 0 1 1570
box -8 -3 32 105
use FILL  FILL_665
timestamp 1681620392
transform 1 0 2872 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_188
timestamp 1681620392
transform -1 0 2896 0 1 1570
box -9 -3 26 105
use FILL  FILL_666
timestamp 1681620392
transform 1 0 2896 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_189
timestamp 1681620392
transform -1 0 2920 0 1 1570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_169
timestamp 1681620392
transform 1 0 2920 0 1 1570
box -8 -3 104 105
use Project_Top_VIA0  Project_Top_VIA0_29
timestamp 1681620392
transform 1 0 3043 0 1 1570
box -10 -3 10 3
use M3_M2  M3_M2_2391
timestamp 1681620392
transform 1 0 132 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2769
timestamp 1681620392
transform 1 0 84 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2392
timestamp 1681620392
transform 1 0 204 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2770
timestamp 1681620392
transform 1 0 180 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2771
timestamp 1681620392
transform 1 0 204 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2772
timestamp 1681620392
transform 1 0 220 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2773
timestamp 1681620392
transform 1 0 228 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2838
timestamp 1681620392
transform 1 0 132 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2839
timestamp 1681620392
transform 1 0 164 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2840
timestamp 1681620392
transform 1 0 172 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2841
timestamp 1681620392
transform 1 0 180 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2842
timestamp 1681620392
transform 1 0 196 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2843
timestamp 1681620392
transform 1 0 212 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2437
timestamp 1681620392
transform 1 0 220 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2393
timestamp 1681620392
transform 1 0 244 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2774
timestamp 1681620392
transform 1 0 244 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2911
timestamp 1681620392
transform 1 0 244 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_2371
timestamp 1681620392
transform 1 0 276 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_2758
timestamp 1681620392
transform 1 0 276 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2844
timestamp 1681620392
transform 1 0 268 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2394
timestamp 1681620392
transform 1 0 284 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2759
timestamp 1681620392
transform 1 0 292 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_2425
timestamp 1681620392
transform 1 0 300 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_2760
timestamp 1681620392
transform 1 0 316 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2775
timestamp 1681620392
transform 1 0 308 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2845
timestamp 1681620392
transform 1 0 300 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2426
timestamp 1681620392
transform 1 0 316 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_2761
timestamp 1681620392
transform 1 0 332 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_2427
timestamp 1681620392
transform 1 0 340 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2351
timestamp 1681620392
transform 1 0 364 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2395
timestamp 1681620392
transform 1 0 364 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2776
timestamp 1681620392
transform 1 0 348 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2846
timestamp 1681620392
transform 1 0 340 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2777
timestamp 1681620392
transform 1 0 372 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2778
timestamp 1681620392
transform 1 0 380 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2847
timestamp 1681620392
transform 1 0 356 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2848
timestamp 1681620392
transform 1 0 364 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2456
timestamp 1681620392
transform 1 0 356 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2457
timestamp 1681620392
transform 1 0 372 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2352
timestamp 1681620392
transform 1 0 396 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2428
timestamp 1681620392
transform 1 0 388 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_2849
timestamp 1681620392
transform 1 0 388 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2762
timestamp 1681620392
transform 1 0 420 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2850
timestamp 1681620392
transform 1 0 420 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2458
timestamp 1681620392
transform 1 0 420 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2372
timestamp 1681620392
transform 1 0 468 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_2779
timestamp 1681620392
transform 1 0 516 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2851
timestamp 1681620392
transform 1 0 468 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2438
timestamp 1681620392
transform 1 0 516 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_2780
timestamp 1681620392
transform 1 0 540 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2396
timestamp 1681620392
transform 1 0 564 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2781
timestamp 1681620392
transform 1 0 556 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2782
timestamp 1681620392
transform 1 0 572 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2852
timestamp 1681620392
transform 1 0 564 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2459
timestamp 1681620392
transform 1 0 564 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_2763
timestamp 1681620392
transform 1 0 588 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2853
timestamp 1681620392
transform 1 0 588 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2373
timestamp 1681620392
transform 1 0 612 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2397
timestamp 1681620392
transform 1 0 620 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2783
timestamp 1681620392
transform 1 0 612 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2439
timestamp 1681620392
transform 1 0 604 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_2764
timestamp 1681620392
transform 1 0 644 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_2460
timestamp 1681620392
transform 1 0 644 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_2784
timestamp 1681620392
transform 1 0 684 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2374
timestamp 1681620392
transform 1 0 716 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2398
timestamp 1681620392
transform 1 0 708 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2785
timestamp 1681620392
transform 1 0 708 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2786
timestamp 1681620392
transform 1 0 716 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2854
timestamp 1681620392
transform 1 0 708 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2855
timestamp 1681620392
transform 1 0 716 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2765
timestamp 1681620392
transform 1 0 740 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_2375
timestamp 1681620392
transform 1 0 764 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_2787
timestamp 1681620392
transform 1 0 764 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2856
timestamp 1681620392
transform 1 0 764 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2857
timestamp 1681620392
transform 1 0 772 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2461
timestamp 1681620392
transform 1 0 764 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2491
timestamp 1681620392
transform 1 0 772 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2399
timestamp 1681620392
transform 1 0 796 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2440
timestamp 1681620392
transform 1 0 788 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_2912
timestamp 1681620392
transform 1 0 788 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2788
timestamp 1681620392
transform 1 0 804 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2462
timestamp 1681620392
transform 1 0 804 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2400
timestamp 1681620392
transform 1 0 852 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2789
timestamp 1681620392
transform 1 0 852 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2441
timestamp 1681620392
transform 1 0 844 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_2858
timestamp 1681620392
transform 1 0 860 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2913
timestamp 1681620392
transform 1 0 836 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2914
timestamp 1681620392
transform 1 0 852 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_2483
timestamp 1681620392
transform 1 0 860 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_2790
timestamp 1681620392
transform 1 0 884 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2442
timestamp 1681620392
transform 1 0 876 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_2915
timestamp 1681620392
transform 1 0 876 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2859
timestamp 1681620392
transform 1 0 892 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2492
timestamp 1681620392
transform 1 0 884 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2401
timestamp 1681620392
transform 1 0 932 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2860
timestamp 1681620392
transform 1 0 908 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2861
timestamp 1681620392
transform 1 0 924 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2791
timestamp 1681620392
transform 1 0 972 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2862
timestamp 1681620392
transform 1 0 948 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2863
timestamp 1681620392
transform 1 0 972 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2916
timestamp 1681620392
transform 1 0 932 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_2463
timestamp 1681620392
transform 1 0 940 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2484
timestamp 1681620392
transform 1 0 932 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_2938
timestamp 1681620392
transform 1 0 940 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_2917
timestamp 1681620392
transform 1 0 964 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_2402
timestamp 1681620392
transform 1 0 988 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2792
timestamp 1681620392
transform 1 0 988 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2864
timestamp 1681620392
transform 1 0 988 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2793
timestamp 1681620392
transform 1 0 1036 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2918
timestamp 1681620392
transform 1 0 1036 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_2493
timestamp 1681620392
transform 1 0 1028 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_2865
timestamp 1681620392
transform 1 0 1044 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2794
timestamp 1681620392
transform 1 0 1076 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2376
timestamp 1681620392
transform 1 0 1132 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_2766
timestamp 1681620392
transform 1 0 1124 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2795
timestamp 1681620392
transform 1 0 1132 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2866
timestamp 1681620392
transform 1 0 1124 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2867
timestamp 1681620392
transform 1 0 1132 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2868
timestamp 1681620392
transform 1 0 1148 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2403
timestamp 1681620392
transform 1 0 1196 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2796
timestamp 1681620392
transform 1 0 1196 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2377
timestamp 1681620392
transform 1 0 1212 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2353
timestamp 1681620392
transform 1 0 1244 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_2797
timestamp 1681620392
transform 1 0 1212 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2429
timestamp 1681620392
transform 1 0 1228 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_2869
timestamp 1681620392
transform 1 0 1220 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2870
timestamp 1681620392
transform 1 0 1228 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2464
timestamp 1681620392
transform 1 0 1204 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_2919
timestamp 1681620392
transform 1 0 1212 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_2430
timestamp 1681620392
transform 1 0 1252 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_2798
timestamp 1681620392
transform 1 0 1260 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2920
timestamp 1681620392
transform 1 0 1236 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2871
timestamp 1681620392
transform 1 0 1276 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2485
timestamp 1681620392
transform 1 0 1268 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2378
timestamp 1681620392
transform 1 0 1292 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2379
timestamp 1681620392
transform 1 0 1308 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_2872
timestamp 1681620392
transform 1 0 1300 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2465
timestamp 1681620392
transform 1 0 1292 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2443
timestamp 1681620392
transform 1 0 1308 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_2873
timestamp 1681620392
transform 1 0 1316 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2799
timestamp 1681620392
transform 1 0 1332 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2466
timestamp 1681620392
transform 1 0 1308 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_2921
timestamp 1681620392
transform 1 0 1316 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_2467
timestamp 1681620392
transform 1 0 1324 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2486
timestamp 1681620392
transform 1 0 1324 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_2922
timestamp 1681620392
transform 1 0 1340 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_2380
timestamp 1681620392
transform 1 0 1372 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2431
timestamp 1681620392
transform 1 0 1364 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2444
timestamp 1681620392
transform 1 0 1356 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_2874
timestamp 1681620392
transform 1 0 1364 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2404
timestamp 1681620392
transform 1 0 1388 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2800
timestamp 1681620392
transform 1 0 1388 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2875
timestamp 1681620392
transform 1 0 1388 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2923
timestamp 1681620392
transform 1 0 1380 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2939
timestamp 1681620392
transform 1 0 1372 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_2494
timestamp 1681620392
transform 1 0 1372 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2468
timestamp 1681620392
transform 1 0 1388 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2432
timestamp 1681620392
transform 1 0 1396 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2495
timestamp 1681620392
transform 1 0 1404 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2354
timestamp 1681620392
transform 1 0 1436 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_2767
timestamp 1681620392
transform 1 0 1428 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2876
timestamp 1681620392
transform 1 0 1428 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2924
timestamp 1681620392
transform 1 0 1436 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_2496
timestamp 1681620392
transform 1 0 1428 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_2877
timestamp 1681620392
transform 1 0 1460 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2445
timestamp 1681620392
transform 1 0 1476 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_2925
timestamp 1681620392
transform 1 0 1476 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2926
timestamp 1681620392
transform 1 0 1484 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2940
timestamp 1681620392
transform 1 0 1468 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_2878
timestamp 1681620392
transform 1 0 1508 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2355
timestamp 1681620392
transform 1 0 1532 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_2801
timestamp 1681620392
transform 1 0 1532 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2802
timestamp 1681620392
transform 1 0 1540 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2503
timestamp 1681620392
transform 1 0 1524 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2497
timestamp 1681620392
transform 1 0 1548 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_2879
timestamp 1681620392
transform 1 0 1564 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2405
timestamp 1681620392
transform 1 0 1604 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2803
timestamp 1681620392
transform 1 0 1604 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2880
timestamp 1681620392
transform 1 0 1588 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2356
timestamp 1681620392
transform 1 0 1628 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2357
timestamp 1681620392
transform 1 0 1644 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2358
timestamp 1681620392
transform 1 0 1724 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2381
timestamp 1681620392
transform 1 0 1668 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2382
timestamp 1681620392
transform 1 0 1692 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2406
timestamp 1681620392
transform 1 0 1660 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2804
timestamp 1681620392
transform 1 0 1620 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2805
timestamp 1681620392
transform 1 0 1708 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2806
timestamp 1681620392
transform 1 0 1724 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2807
timestamp 1681620392
transform 1 0 1740 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2881
timestamp 1681620392
transform 1 0 1612 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2882
timestamp 1681620392
transform 1 0 1620 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2883
timestamp 1681620392
transform 1 0 1660 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2469
timestamp 1681620392
transform 1 0 1588 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_2927
timestamp 1681620392
transform 1 0 1604 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_2470
timestamp 1681620392
transform 1 0 1612 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2487
timestamp 1681620392
transform 1 0 1604 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2446
timestamp 1681620392
transform 1 0 1684 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2504
timestamp 1681620392
transform 1 0 1700 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2359
timestamp 1681620392
transform 1 0 1772 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2407
timestamp 1681620392
transform 1 0 1764 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2408
timestamp 1681620392
transform 1 0 1804 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2808
timestamp 1681620392
transform 1 0 1764 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2809
timestamp 1681620392
transform 1 0 1852 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2447
timestamp 1681620392
transform 1 0 1764 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2409
timestamp 1681620392
transform 1 0 1908 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2360
timestamp 1681620392
transform 1 0 1940 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2383
timestamp 1681620392
transform 1 0 1940 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2410
timestamp 1681620392
transform 1 0 1948 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2810
timestamp 1681620392
transform 1 0 1884 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2811
timestamp 1681620392
transform 1 0 1908 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2812
timestamp 1681620392
transform 1 0 1932 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2884
timestamp 1681620392
transform 1 0 1772 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2885
timestamp 1681620392
transform 1 0 1804 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2886
timestamp 1681620392
transform 1 0 1868 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2928
timestamp 1681620392
transform 1 0 1764 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_2505
timestamp 1681620392
transform 1 0 1780 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2506
timestamp 1681620392
transform 1 0 1836 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2433
timestamp 1681620392
transform 1 0 1940 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_2813
timestamp 1681620392
transform 1 0 1956 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2361
timestamp 1681620392
transform 1 0 2020 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2411
timestamp 1681620392
transform 1 0 1996 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2814
timestamp 1681620392
transform 1 0 1980 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2815
timestamp 1681620392
transform 1 0 1996 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2887
timestamp 1681620392
transform 1 0 1892 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2888
timestamp 1681620392
transform 1 0 1916 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2889
timestamp 1681620392
transform 1 0 1940 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2890
timestamp 1681620392
transform 1 0 1964 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2471
timestamp 1681620392
transform 1 0 1908 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2448
timestamp 1681620392
transform 1 0 1980 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2362
timestamp 1681620392
transform 1 0 2092 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2412
timestamp 1681620392
transform 1 0 2092 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2413
timestamp 1681620392
transform 1 0 2140 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2816
timestamp 1681620392
transform 1 0 2092 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2891
timestamp 1681620392
transform 1 0 2036 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2892
timestamp 1681620392
transform 1 0 2076 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2893
timestamp 1681620392
transform 1 0 2132 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2472
timestamp 1681620392
transform 1 0 1940 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2473
timestamp 1681620392
transform 1 0 1964 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2488
timestamp 1681620392
transform 1 0 1972 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2507
timestamp 1681620392
transform 1 0 2156 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2434
timestamp 1681620392
transform 1 0 2196 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2363
timestamp 1681620392
transform 1 0 2220 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2384
timestamp 1681620392
transform 1 0 2212 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2414
timestamp 1681620392
transform 1 0 2220 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2817
timestamp 1681620392
transform 1 0 2212 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2818
timestamp 1681620392
transform 1 0 2220 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2894
timestamp 1681620392
transform 1 0 2188 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2895
timestamp 1681620392
transform 1 0 2204 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2896
timestamp 1681620392
transform 1 0 2212 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2474
timestamp 1681620392
transform 1 0 2188 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_2929
timestamp 1681620392
transform 1 0 2196 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_2475
timestamp 1681620392
transform 1 0 2212 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2498
timestamp 1681620392
transform 1 0 2204 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2508
timestamp 1681620392
transform 1 0 2212 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2385
timestamp 1681620392
transform 1 0 2260 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2415
timestamp 1681620392
transform 1 0 2252 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2819
timestamp 1681620392
transform 1 0 2252 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2449
timestamp 1681620392
transform 1 0 2252 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_2930
timestamp 1681620392
transform 1 0 2252 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2820
timestamp 1681620392
transform 1 0 2276 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2476
timestamp 1681620392
transform 1 0 2276 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2364
timestamp 1681620392
transform 1 0 2292 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2416
timestamp 1681620392
transform 1 0 2316 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2821
timestamp 1681620392
transform 1 0 2292 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2822
timestamp 1681620392
transform 1 0 2380 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2897
timestamp 1681620392
transform 1 0 2316 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2450
timestamp 1681620392
transform 1 0 2340 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_2898
timestamp 1681620392
transform 1 0 2372 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2451
timestamp 1681620392
transform 1 0 2380 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2386
timestamp 1681620392
transform 1 0 2412 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_2823
timestamp 1681620392
transform 1 0 2404 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2452
timestamp 1681620392
transform 1 0 2404 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2477
timestamp 1681620392
transform 1 0 2372 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_2931
timestamp 1681620392
transform 1 0 2380 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_2478
timestamp 1681620392
transform 1 0 2388 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_2932
timestamp 1681620392
transform 1 0 2412 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_2499
timestamp 1681620392
transform 1 0 2372 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2387
timestamp 1681620392
transform 1 0 2436 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2417
timestamp 1681620392
transform 1 0 2428 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2824
timestamp 1681620392
transform 1 0 2428 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2825
timestamp 1681620392
transform 1 0 2436 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2899
timestamp 1681620392
transform 1 0 2436 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2418
timestamp 1681620392
transform 1 0 2452 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2826
timestamp 1681620392
transform 1 0 2452 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2453
timestamp 1681620392
transform 1 0 2452 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_2933
timestamp 1681620392
transform 1 0 2452 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_2500
timestamp 1681620392
transform 1 0 2444 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2479
timestamp 1681620392
transform 1 0 2460 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2365
timestamp 1681620392
transform 1 0 2580 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2388
timestamp 1681620392
transform 1 0 2500 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2419
timestamp 1681620392
transform 1 0 2500 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2827
timestamp 1681620392
transform 1 0 2580 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2900
timestamp 1681620392
transform 1 0 2484 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2901
timestamp 1681620392
transform 1 0 2500 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2902
timestamp 1681620392
transform 1 0 2556 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2509
timestamp 1681620392
transform 1 0 2564 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_2828
timestamp 1681620392
transform 1 0 2604 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2510
timestamp 1681620392
transform 1 0 2604 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_2829
timestamp 1681620392
transform 1 0 2620 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2903
timestamp 1681620392
transform 1 0 2620 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2366
timestamp 1681620392
transform 1 0 2724 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2389
timestamp 1681620392
transform 1 0 2708 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2420
timestamp 1681620392
transform 1 0 2644 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2367
timestamp 1681620392
transform 1 0 2756 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2421
timestamp 1681620392
transform 1 0 2740 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2435
timestamp 1681620392
transform 1 0 2700 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_2830
timestamp 1681620392
transform 1 0 2724 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2831
timestamp 1681620392
transform 1 0 2740 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2832
timestamp 1681620392
transform 1 0 2756 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2904
timestamp 1681620392
transform 1 0 2636 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2905
timestamp 1681620392
transform 1 0 2644 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2906
timestamp 1681620392
transform 1 0 2700 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2436
timestamp 1681620392
transform 1 0 2772 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_2768
timestamp 1681620392
transform 1 0 2788 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2833
timestamp 1681620392
transform 1 0 2780 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2834
timestamp 1681620392
transform 1 0 2796 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2454
timestamp 1681620392
transform 1 0 2780 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2455
timestamp 1681620392
transform 1 0 2812 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_2934
timestamp 1681620392
transform 1 0 2780 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_2511
timestamp 1681620392
transform 1 0 2764 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2480
timestamp 1681620392
transform 1 0 2796 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2489
timestamp 1681620392
transform 1 0 2804 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2512
timestamp 1681620392
transform 1 0 2796 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2368
timestamp 1681620392
transform 1 0 2836 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2422
timestamp 1681620392
transform 1 0 2836 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2835
timestamp 1681620392
transform 1 0 2836 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_2390
timestamp 1681620392
transform 1 0 2852 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2369
timestamp 1681620392
transform 1 0 2884 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2423
timestamp 1681620392
transform 1 0 2868 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2836
timestamp 1681620392
transform 1 0 2868 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2907
timestamp 1681620392
transform 1 0 2844 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2908
timestamp 1681620392
transform 1 0 2860 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2424
timestamp 1681620392
transform 1 0 2900 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2909
timestamp 1681620392
transform 1 0 2892 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2935
timestamp 1681620392
transform 1 0 2868 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_2481
timestamp 1681620392
transform 1 0 2892 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_2936
timestamp 1681620392
transform 1 0 2900 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_2490
timestamp 1681620392
transform 1 0 2868 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_2941
timestamp 1681620392
transform 1 0 2884 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_2501
timestamp 1681620392
transform 1 0 2852 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2502
timestamp 1681620392
transform 1 0 2892 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_2910
timestamp 1681620392
transform 1 0 2916 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_2482
timestamp 1681620392
transform 1 0 2916 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2370
timestamp 1681620392
transform 1 0 2932 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_2837
timestamp 1681620392
transform 1 0 2940 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2937
timestamp 1681620392
transform 1 0 2956 0 1 1515
box -2 -2 2 2
use Project_Top_VIA0  Project_Top_VIA0_30
timestamp 1681620392
transform 1 0 24 0 1 1470
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_162
timestamp 1681620392
transform 1 0 72 0 -1 1570
box -8 -3 104 105
use INVX2  INVX2_176
timestamp 1681620392
transform -1 0 184 0 -1 1570
box -9 -3 26 105
use OAI22X1  OAI22X1_41
timestamp 1681620392
transform 1 0 184 0 -1 1570
box -8 -3 46 105
use NAND2X1  NAND2X1_145
timestamp 1681620392
transform 1 0 224 0 -1 1570
box -8 -3 32 105
use FILL  FILL_562
timestamp 1681620392
transform 1 0 248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_563
timestamp 1681620392
transform 1 0 256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_564
timestamp 1681620392
transform 1 0 264 0 -1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_52
timestamp 1681620392
transform 1 0 272 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_53
timestamp 1681620392
transform 1 0 296 0 -1 1570
box -8 -3 32 105
use FILL  FILL_565
timestamp 1681620392
transform 1 0 320 0 -1 1570
box -8 -3 16 105
use FILL  FILL_566
timestamp 1681620392
transform 1 0 328 0 -1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_54
timestamp 1681620392
transform 1 0 336 0 -1 1570
box -8 -3 32 105
use INVX2  INVX2_177
timestamp 1681620392
transform -1 0 376 0 -1 1570
box -9 -3 26 105
use FILL  FILL_567
timestamp 1681620392
transform 1 0 376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_568
timestamp 1681620392
transform 1 0 384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_569
timestamp 1681620392
transform 1 0 392 0 -1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_55
timestamp 1681620392
transform -1 0 424 0 -1 1570
box -8 -3 32 105
use FILL  FILL_570
timestamp 1681620392
transform 1 0 424 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_163
timestamp 1681620392
transform -1 0 528 0 -1 1570
box -8 -3 104 105
use FILL  FILL_571
timestamp 1681620392
transform 1 0 528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_572
timestamp 1681620392
transform 1 0 536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_573
timestamp 1681620392
transform 1 0 544 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_178
timestamp 1681620392
transform 1 0 552 0 -1 1570
box -9 -3 26 105
use NOR2X1  NOR2X1_56
timestamp 1681620392
transform -1 0 592 0 -1 1570
box -8 -3 32 105
use FILL  FILL_574
timestamp 1681620392
transform 1 0 592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_575
timestamp 1681620392
transform 1 0 600 0 -1 1570
box -8 -3 16 105
use FILL  FILL_576
timestamp 1681620392
transform 1 0 608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_577
timestamp 1681620392
transform 1 0 616 0 -1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_57
timestamp 1681620392
transform -1 0 648 0 -1 1570
box -8 -3 32 105
use FILL  FILL_578
timestamp 1681620392
transform 1 0 648 0 -1 1570
box -8 -3 16 105
use FILL  FILL_579
timestamp 1681620392
transform 1 0 656 0 -1 1570
box -8 -3 16 105
use FILL  FILL_581
timestamp 1681620392
transform 1 0 664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_584
timestamp 1681620392
transform 1 0 672 0 -1 1570
box -8 -3 16 105
use FILL  FILL_585
timestamp 1681620392
transform 1 0 680 0 -1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_147
timestamp 1681620392
transform -1 0 712 0 -1 1570
box -8 -3 32 105
use AOI21X1  AOI21X1_14
timestamp 1681620392
transform 1 0 712 0 -1 1570
box -7 -3 39 105
use FILL  FILL_586
timestamp 1681620392
transform 1 0 744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_587
timestamp 1681620392
transform 1 0 752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_589
timestamp 1681620392
transform 1 0 760 0 -1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_149
timestamp 1681620392
transform 1 0 768 0 -1 1570
box -8 -3 32 105
use FILL  FILL_592
timestamp 1681620392
transform 1 0 792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_593
timestamp 1681620392
transform 1 0 800 0 -1 1570
box -8 -3 16 105
use FILL  FILL_595
timestamp 1681620392
transform 1 0 808 0 -1 1570
box -8 -3 16 105
use FILL  FILL_597
timestamp 1681620392
transform 1 0 816 0 -1 1570
box -8 -3 16 105
use FILL  FILL_601
timestamp 1681620392
transform 1 0 824 0 -1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_152
timestamp 1681620392
transform 1 0 832 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_153
timestamp 1681620392
transform 1 0 856 0 -1 1570
box -8 -3 32 105
use FILL  FILL_602
timestamp 1681620392
transform 1 0 880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_603
timestamp 1681620392
transform 1 0 888 0 -1 1570
box -8 -3 16 105
use AND2X2  AND2X2_14
timestamp 1681620392
transform 1 0 896 0 -1 1570
box -8 -3 40 105
use FILL  FILL_604
timestamp 1681620392
transform 1 0 928 0 -1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_56
timestamp 1681620392
transform 1 0 936 0 -1 1570
box -8 -3 40 105
use INVX2  INVX2_181
timestamp 1681620392
transform 1 0 968 0 -1 1570
box -9 -3 26 105
use FILL  FILL_605
timestamp 1681620392
transform 1 0 984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_606
timestamp 1681620392
transform 1 0 992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_607
timestamp 1681620392
transform 1 0 1000 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_167
timestamp 1681620392
transform 1 0 1008 0 -1 1570
box -8 -3 34 105
use FILL  FILL_608
timestamp 1681620392
transform 1 0 1040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_609
timestamp 1681620392
transform 1 0 1048 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_182
timestamp 1681620392
transform -1 0 1072 0 -1 1570
box -9 -3 26 105
use FILL  FILL_610
timestamp 1681620392
transform 1 0 1072 0 -1 1570
box -8 -3 16 105
use FILL  FILL_611
timestamp 1681620392
transform 1 0 1080 0 -1 1570
box -8 -3 16 105
use FILL  FILL_612
timestamp 1681620392
transform 1 0 1088 0 -1 1570
box -8 -3 16 105
use FILL  FILL_613
timestamp 1681620392
transform 1 0 1096 0 -1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_60
timestamp 1681620392
transform 1 0 1104 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_61
timestamp 1681620392
transform 1 0 1128 0 -1 1570
box -8 -3 32 105
use FILL  FILL_614
timestamp 1681620392
transform 1 0 1152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_615
timestamp 1681620392
transform 1 0 1160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_616
timestamp 1681620392
transform 1 0 1168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_617
timestamp 1681620392
transform 1 0 1176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_618
timestamp 1681620392
transform 1 0 1184 0 -1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_154
timestamp 1681620392
transform 1 0 1192 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_156
timestamp 1681620392
transform 1 0 1216 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_157
timestamp 1681620392
transform -1 0 1264 0 -1 1570
box -8 -3 32 105
use FILL  FILL_623
timestamp 1681620392
transform 1 0 1264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_627
timestamp 1681620392
transform 1 0 1272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_628
timestamp 1681620392
transform 1 0 1280 0 -1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_161
timestamp 1681620392
transform 1 0 1288 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_162
timestamp 1681620392
transform -1 0 1336 0 -1 1570
box -8 -3 32 105
use FILL  FILL_629
timestamp 1681620392
transform 1 0 1336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_630
timestamp 1681620392
transform 1 0 1344 0 -1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_58
timestamp 1681620392
transform 1 0 1352 0 -1 1570
box -8 -3 40 105
use FILL  FILL_631
timestamp 1681620392
transform 1 0 1384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_632
timestamp 1681620392
transform 1 0 1392 0 -1 1570
box -8 -3 16 105
use AOI21X1  AOI21X1_16
timestamp 1681620392
transform 1 0 1400 0 -1 1570
box -7 -3 39 105
use FILL  FILL_633
timestamp 1681620392
transform 1 0 1432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_634
timestamp 1681620392
transform 1 0 1440 0 -1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_59
timestamp 1681620392
transform 1 0 1448 0 -1 1570
box -8 -3 40 105
use FILL  FILL_638
timestamp 1681620392
transform 1 0 1480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_640
timestamp 1681620392
transform 1 0 1488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_642
timestamp 1681620392
transform 1 0 1496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_667
timestamp 1681620392
transform 1 0 1504 0 -1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_167
timestamp 1681620392
transform -1 0 1536 0 -1 1570
box -8 -3 32 105
use FILL  FILL_668
timestamp 1681620392
transform 1 0 1536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_669
timestamp 1681620392
transform 1 0 1544 0 -1 1570
box -8 -3 16 105
use FILL  FILL_670
timestamp 1681620392
transform 1 0 1552 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_190
timestamp 1681620392
transform 1 0 1560 0 -1 1570
box -9 -3 26 105
use OAI21X1  OAI21X1_173
timestamp 1681620392
transform 1 0 1576 0 -1 1570
box -8 -3 34 105
use INVX2  INVX2_191
timestamp 1681620392
transform -1 0 1624 0 -1 1570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_170
timestamp 1681620392
transform -1 0 1720 0 -1 1570
box -8 -3 104 105
use INVX2  INVX2_192
timestamp 1681620392
transform 1 0 1720 0 -1 1570
box -9 -3 26 105
use OAI21X1  OAI21X1_174
timestamp 1681620392
transform 1 0 1736 0 -1 1570
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_171
timestamp 1681620392
transform -1 0 1864 0 -1 1570
box -8 -3 104 105
use BUFX2  BUFX2_25
timestamp 1681620392
transform 1 0 1864 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_26
timestamp 1681620392
transform 1 0 1888 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_27
timestamp 1681620392
transform 1 0 1912 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_28
timestamp 1681620392
transform 1 0 1936 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_29
timestamp 1681620392
transform 1 0 1960 0 -1 1570
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_172
timestamp 1681620392
transform 1 0 1984 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_173
timestamp 1681620392
transform 1 0 2080 0 -1 1570
box -8 -3 104 105
use INVX2  INVX2_193
timestamp 1681620392
transform 1 0 2176 0 -1 1570
box -9 -3 26 105
use NAND2X1  NAND2X1_168
timestamp 1681620392
transform -1 0 2216 0 -1 1570
box -8 -3 32 105
use OAI21X1  OAI21X1_175
timestamp 1681620392
transform 1 0 2216 0 -1 1570
box -8 -3 34 105
use NAND2X1  NAND2X1_169
timestamp 1681620392
transform -1 0 2272 0 -1 1570
box -8 -3 32 105
use FILL  FILL_671
timestamp 1681620392
transform 1 0 2272 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_174
timestamp 1681620392
transform 1 0 2280 0 -1 1570
box -8 -3 104 105
use OAI21X1  OAI21X1_176
timestamp 1681620392
transform -1 0 2408 0 -1 1570
box -8 -3 34 105
use NAND2X1  NAND2X1_170
timestamp 1681620392
transform -1 0 2432 0 -1 1570
box -8 -3 32 105
use M3_M2  M3_M2_2513
timestamp 1681620392
transform 1 0 2452 0 1 1475
box -3 -3 3 3
use NAND2X1  NAND2X1_171
timestamp 1681620392
transform 1 0 2432 0 -1 1570
box -8 -3 32 105
use FILL  FILL_672
timestamp 1681620392
transform 1 0 2456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_673
timestamp 1681620392
transform 1 0 2464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_674
timestamp 1681620392
transform 1 0 2472 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_2514
timestamp 1681620392
transform 1 0 2508 0 1 1475
box -3 -3 3 3
use INVX2  INVX2_194
timestamp 1681620392
transform 1 0 2480 0 -1 1570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_175
timestamp 1681620392
transform -1 0 2592 0 -1 1570
box -8 -3 104 105
use FILL  FILL_675
timestamp 1681620392
transform 1 0 2592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_676
timestamp 1681620392
transform 1 0 2600 0 -1 1570
box -8 -3 16 105
use FILL  FILL_677
timestamp 1681620392
transform 1 0 2608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_678
timestamp 1681620392
transform 1 0 2616 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_2515
timestamp 1681620392
transform 1 0 2636 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2516
timestamp 1681620392
transform 1 0 2692 0 1 1475
box -3 -3 3 3
use INVX2  INVX2_195
timestamp 1681620392
transform 1 0 2624 0 -1 1570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_176
timestamp 1681620392
transform -1 0 2736 0 -1 1570
box -8 -3 104 105
use M3_M2  M3_M2_2517
timestamp 1681620392
transform 1 0 2764 0 1 1475
box -3 -3 3 3
use INVX2  INVX2_196
timestamp 1681620392
transform 1 0 2736 0 -1 1570
box -9 -3 26 105
use OAI21X1  OAI21X1_177
timestamp 1681620392
transform 1 0 2752 0 -1 1570
box -8 -3 34 105
use NOR2X1  NOR2X1_65
timestamp 1681620392
transform 1 0 2784 0 -1 1570
box -8 -3 32 105
use INVX2  INVX2_197
timestamp 1681620392
transform -1 0 2824 0 -1 1570
box -9 -3 26 105
use FILL  FILL_679
timestamp 1681620392
transform 1 0 2824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_680
timestamp 1681620392
transform 1 0 2832 0 -1 1570
box -8 -3 16 105
use AND2X2  AND2X2_15
timestamp 1681620392
transform -1 0 2872 0 -1 1570
box -8 -3 40 105
use M3_M2  M3_M2_2518
timestamp 1681620392
transform 1 0 2884 0 1 1475
box -3 -3 3 3
use NAND3X1  NAND3X1_63
timestamp 1681620392
transform -1 0 2904 0 -1 1570
box -8 -3 40 105
use FILL  FILL_681
timestamp 1681620392
transform 1 0 2904 0 -1 1570
box -8 -3 16 105
use FILL  FILL_682
timestamp 1681620392
transform 1 0 2912 0 -1 1570
box -8 -3 16 105
use FILL  FILL_683
timestamp 1681620392
transform 1 0 2920 0 -1 1570
box -8 -3 16 105
use FILL  FILL_684
timestamp 1681620392
transform 1 0 2928 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_2519
timestamp 1681620392
transform 1 0 2964 0 1 1475
box -3 -3 3 3
use NAND2X1  NAND2X1_172
timestamp 1681620392
transform 1 0 2936 0 -1 1570
box -8 -3 32 105
use FILL  FILL_685
timestamp 1681620392
transform 1 0 2960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_686
timestamp 1681620392
transform 1 0 2968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_687
timestamp 1681620392
transform 1 0 2976 0 -1 1570
box -8 -3 16 105
use FILL  FILL_688
timestamp 1681620392
transform 1 0 2984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_689
timestamp 1681620392
transform 1 0 2992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_690
timestamp 1681620392
transform 1 0 3000 0 -1 1570
box -8 -3 16 105
use FILL  FILL_691
timestamp 1681620392
transform 1 0 3008 0 -1 1570
box -8 -3 16 105
use Project_Top_VIA0  Project_Top_VIA0_31
timestamp 1681620392
transform 1 0 3067 0 1 1470
box -10 -3 10 3
use M2_M1  M2_M1_3060
timestamp 1681620392
transform 1 0 92 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3134
timestamp 1681620392
transform 1 0 140 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_2552
timestamp 1681620392
transform 1 0 164 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_2983
timestamp 1681620392
transform 1 0 164 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2984
timestamp 1681620392
transform 1 0 172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3135
timestamp 1681620392
transform 1 0 180 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_2553
timestamp 1681620392
transform 1 0 196 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_2985
timestamp 1681620392
transform 1 0 196 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2986
timestamp 1681620392
transform 1 0 204 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2946
timestamp 1681620392
transform 1 0 220 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_2572
timestamp 1681620392
transform 1 0 228 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_3061
timestamp 1681620392
transform 1 0 228 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2947
timestamp 1681620392
transform 1 0 244 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_2573
timestamp 1681620392
transform 1 0 244 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_3062
timestamp 1681620392
transform 1 0 252 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2987
timestamp 1681620392
transform 1 0 276 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2948
timestamp 1681620392
transform 1 0 292 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_2574
timestamp 1681620392
transform 1 0 292 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_3063
timestamp 1681620392
transform 1 0 292 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2592
timestamp 1681620392
transform 1 0 308 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2535
timestamp 1681620392
transform 1 0 332 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_2988
timestamp 1681620392
transform 1 0 332 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3064
timestamp 1681620392
transform 1 0 316 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2611
timestamp 1681620392
transform 1 0 292 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2593
timestamp 1681620392
transform 1 0 324 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_3065
timestamp 1681620392
transform 1 0 332 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2639
timestamp 1681620392
transform 1 0 324 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_2949
timestamp 1681620392
transform 1 0 348 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2989
timestamp 1681620392
transform 1 0 356 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3066
timestamp 1681620392
transform 1 0 356 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2612
timestamp 1681620392
transform 1 0 348 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2640
timestamp 1681620392
transform 1 0 356 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_2950
timestamp 1681620392
transform 1 0 372 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_2575
timestamp 1681620392
transform 1 0 372 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_2990
timestamp 1681620392
transform 1 0 396 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2991
timestamp 1681620392
transform 1 0 404 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2942
timestamp 1681620392
transform 1 0 420 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_3067
timestamp 1681620392
transform 1 0 412 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2536
timestamp 1681620392
transform 1 0 428 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_2951
timestamp 1681620392
transform 1 0 428 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_2576
timestamp 1681620392
transform 1 0 428 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_2992
timestamp 1681620392
transform 1 0 436 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_2613
timestamp 1681620392
transform 1 0 428 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2537
timestamp 1681620392
transform 1 0 476 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_2952
timestamp 1681620392
transform 1 0 508 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3068
timestamp 1681620392
transform 1 0 500 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2953
timestamp 1681620392
transform 1 0 532 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3069
timestamp 1681620392
transform 1 0 524 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2993
timestamp 1681620392
transform 1 0 540 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_2520
timestamp 1681620392
transform 1 0 668 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_2994
timestamp 1681620392
transform 1 0 556 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2995
timestamp 1681620392
transform 1 0 572 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2996
timestamp 1681620392
transform 1 0 588 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2997
timestamp 1681620392
transform 1 0 620 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3070
timestamp 1681620392
transform 1 0 564 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2594
timestamp 1681620392
transform 1 0 572 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_3071
timestamp 1681620392
transform 1 0 580 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3072
timestamp 1681620392
transform 1 0 668 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2614
timestamp 1681620392
transform 1 0 580 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2521
timestamp 1681620392
transform 1 0 700 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2526
timestamp 1681620392
transform 1 0 716 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_2943
timestamp 1681620392
transform 1 0 700 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_2954
timestamp 1681620392
transform 1 0 692 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2955
timestamp 1681620392
transform 1 0 716 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2998
timestamp 1681620392
transform 1 0 708 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2999
timestamp 1681620392
transform 1 0 724 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3000
timestamp 1681620392
transform 1 0 732 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3001
timestamp 1681620392
transform 1 0 740 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_2595
timestamp 1681620392
transform 1 0 700 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2615
timestamp 1681620392
transform 1 0 692 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2616
timestamp 1681620392
transform 1 0 724 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2538
timestamp 1681620392
transform 1 0 772 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_2956
timestamp 1681620392
transform 1 0 772 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2957
timestamp 1681620392
transform 1 0 780 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3073
timestamp 1681620392
transform 1 0 756 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2596
timestamp 1681620392
transform 1 0 764 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2641
timestamp 1681620392
transform 1 0 756 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2597
timestamp 1681620392
transform 1 0 788 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2554
timestamp 1681620392
transform 1 0 812 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_3002
timestamp 1681620392
transform 1 0 812 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3074
timestamp 1681620392
transform 1 0 796 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3075
timestamp 1681620392
transform 1 0 804 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2617
timestamp 1681620392
transform 1 0 804 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2527
timestamp 1681620392
transform 1 0 828 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2539
timestamp 1681620392
transform 1 0 860 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_2958
timestamp 1681620392
transform 1 0 828 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_2555
timestamp 1681620392
transform 1 0 844 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_2959
timestamp 1681620392
transform 1 0 860 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3003
timestamp 1681620392
transform 1 0 844 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_2528
timestamp 1681620392
transform 1 0 892 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_2960
timestamp 1681620392
transform 1 0 892 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3004
timestamp 1681620392
transform 1 0 884 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3076
timestamp 1681620392
transform 1 0 860 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3077
timestamp 1681620392
transform 1 0 892 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2618
timestamp 1681620392
transform 1 0 884 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2529
timestamp 1681620392
transform 1 0 948 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_2944
timestamp 1681620392
transform 1 0 932 0 1 1435
box -2 -2 2 2
use M3_M2  M3_M2_2556
timestamp 1681620392
transform 1 0 932 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_2961
timestamp 1681620392
transform 1 0 940 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2962
timestamp 1681620392
transform 1 0 948 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3005
timestamp 1681620392
transform 1 0 924 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_2557
timestamp 1681620392
transform 1 0 964 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_3078
timestamp 1681620392
transform 1 0 964 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3079
timestamp 1681620392
transform 1 0 972 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2540
timestamp 1681620392
transform 1 0 1004 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_2963
timestamp 1681620392
transform 1 0 1004 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_2577
timestamp 1681620392
transform 1 0 988 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2598
timestamp 1681620392
transform 1 0 996 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2642
timestamp 1681620392
transform 1 0 988 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_3006
timestamp 1681620392
transform 1 0 1028 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_2578
timestamp 1681620392
transform 1 0 1036 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2558
timestamp 1681620392
transform 1 0 1140 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_3007
timestamp 1681620392
transform 1 0 1100 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3008
timestamp 1681620392
transform 1 0 1132 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3009
timestamp 1681620392
transform 1 0 1140 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3080
timestamp 1681620392
transform 1 0 1012 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3081
timestamp 1681620392
transform 1 0 1036 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3082
timestamp 1681620392
transform 1 0 1052 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3083
timestamp 1681620392
transform 1 0 1140 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2559
timestamp 1681620392
transform 1 0 1164 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_3010
timestamp 1681620392
transform 1 0 1156 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_2522
timestamp 1681620392
transform 1 0 1188 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2560
timestamp 1681620392
transform 1 0 1204 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2561
timestamp 1681620392
transform 1 0 1236 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_3011
timestamp 1681620392
transform 1 0 1204 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3012
timestamp 1681620392
transform 1 0 1220 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3013
timestamp 1681620392
transform 1 0 1236 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3084
timestamp 1681620392
transform 1 0 1188 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3085
timestamp 1681620392
transform 1 0 1196 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2599
timestamp 1681620392
transform 1 0 1204 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_3086
timestamp 1681620392
transform 1 0 1228 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2619
timestamp 1681620392
transform 1 0 1196 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2620
timestamp 1681620392
transform 1 0 1228 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2541
timestamp 1681620392
transform 1 0 1276 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_2964
timestamp 1681620392
transform 1 0 1276 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_2542
timestamp 1681620392
transform 1 0 1316 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_2945
timestamp 1681620392
transform 1 0 1324 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_2965
timestamp 1681620392
transform 1 0 1300 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2966
timestamp 1681620392
transform 1 0 1308 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_2562
timestamp 1681620392
transform 1 0 1324 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_2967
timestamp 1681620392
transform 1 0 1332 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_2563
timestamp 1681620392
transform 1 0 1340 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_3014
timestamp 1681620392
transform 1 0 1284 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_2579
timestamp 1681620392
transform 1 0 1300 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_3015
timestamp 1681620392
transform 1 0 1316 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_2600
timestamp 1681620392
transform 1 0 1300 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_3016
timestamp 1681620392
transform 1 0 1348 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_2580
timestamp 1681620392
transform 1 0 1356 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_2968
timestamp 1681620392
transform 1 0 1380 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3017
timestamp 1681620392
transform 1 0 1364 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3087
timestamp 1681620392
transform 1 0 1340 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2601
timestamp 1681620392
transform 1 0 1348 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_3088
timestamp 1681620392
transform 1 0 1356 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2643
timestamp 1681620392
transform 1 0 1340 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2621
timestamp 1681620392
transform 1 0 1372 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_2969
timestamp 1681620392
transform 1 0 1388 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3089
timestamp 1681620392
transform 1 0 1388 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2644
timestamp 1681620392
transform 1 0 1396 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_2970
timestamp 1681620392
transform 1 0 1420 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_2543
timestamp 1681620392
transform 1 0 1436 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_3018
timestamp 1681620392
transform 1 0 1452 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3090
timestamp 1681620392
transform 1 0 1444 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2523
timestamp 1681620392
transform 1 0 1484 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2544
timestamp 1681620392
transform 1 0 1476 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_2971
timestamp 1681620392
transform 1 0 1476 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_2524
timestamp 1681620392
transform 1 0 1716 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_3019
timestamp 1681620392
transform 1 0 1476 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3020
timestamp 1681620392
transform 1 0 1492 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3021
timestamp 1681620392
transform 1 0 1508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3022
timestamp 1681620392
transform 1 0 1524 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3023
timestamp 1681620392
transform 1 0 1556 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3024
timestamp 1681620392
transform 1 0 1620 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3025
timestamp 1681620392
transform 1 0 1676 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3026
timestamp 1681620392
transform 1 0 1716 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3091
timestamp 1681620392
transform 1 0 1476 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3092
timestamp 1681620392
transform 1 0 1500 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3093
timestamp 1681620392
transform 1 0 1516 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3094
timestamp 1681620392
transform 1 0 1604 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2622
timestamp 1681620392
transform 1 0 1500 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2602
timestamp 1681620392
transform 1 0 1620 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2603
timestamp 1681620392
transform 1 0 1652 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_3095
timestamp 1681620392
transform 1 0 1700 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2623
timestamp 1681620392
transform 1 0 1556 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2624
timestamp 1681620392
transform 1 0 1700 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_3027
timestamp 1681620392
transform 1 0 1740 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3028
timestamp 1681620392
transform 1 0 1764 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3096
timestamp 1681620392
transform 1 0 1732 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3097
timestamp 1681620392
transform 1 0 1756 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2525
timestamp 1681620392
transform 1 0 1868 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_3029
timestamp 1681620392
transform 1 0 1844 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3098
timestamp 1681620392
transform 1 0 1780 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3099
timestamp 1681620392
transform 1 0 1796 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2604
timestamp 1681620392
transform 1 0 1868 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2625
timestamp 1681620392
transform 1 0 1780 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2626
timestamp 1681620392
transform 1 0 1812 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2645
timestamp 1681620392
transform 1 0 1796 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_3030
timestamp 1681620392
transform 1 0 1892 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_2605
timestamp 1681620392
transform 1 0 1892 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_3100
timestamp 1681620392
transform 1 0 1908 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2530
timestamp 1681620392
transform 1 0 1956 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2531
timestamp 1681620392
transform 1 0 2036 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2545
timestamp 1681620392
transform 1 0 1956 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_2972
timestamp 1681620392
transform 1 0 1956 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3031
timestamp 1681620392
transform 1 0 1996 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3101
timestamp 1681620392
transform 1 0 1956 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3102
timestamp 1681620392
transform 1 0 1972 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2627
timestamp 1681620392
transform 1 0 1956 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2628
timestamp 1681620392
transform 1 0 1996 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2646
timestamp 1681620392
transform 1 0 1948 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2546
timestamp 1681620392
transform 1 0 2076 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2547
timestamp 1681620392
transform 1 0 2116 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_2973
timestamp 1681620392
transform 1 0 2084 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_2564
timestamp 1681620392
transform 1 0 2100 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_3032
timestamp 1681620392
transform 1 0 2068 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3033
timestamp 1681620392
transform 1 0 2076 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3103
timestamp 1681620392
transform 1 0 2068 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2629
timestamp 1681620392
transform 1 0 2068 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2581
timestamp 1681620392
transform 1 0 2084 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2565
timestamp 1681620392
transform 1 0 2132 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_2974
timestamp 1681620392
transform 1 0 2140 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3034
timestamp 1681620392
transform 1 0 2100 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3035
timestamp 1681620392
transform 1 0 2116 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_2582
timestamp 1681620392
transform 1 0 2124 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_3036
timestamp 1681620392
transform 1 0 2132 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3104
timestamp 1681620392
transform 1 0 2084 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3105
timestamp 1681620392
transform 1 0 2108 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2606
timestamp 1681620392
transform 1 0 2116 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_3106
timestamp 1681620392
transform 1 0 2124 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3107
timestamp 1681620392
transform 1 0 2132 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2630
timestamp 1681620392
transform 1 0 2108 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2647
timestamp 1681620392
transform 1 0 2172 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2532
timestamp 1681620392
transform 1 0 2204 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_2975
timestamp 1681620392
transform 1 0 2196 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_2548
timestamp 1681620392
transform 1 0 2316 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_2976
timestamp 1681620392
transform 1 0 2316 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3037
timestamp 1681620392
transform 1 0 2204 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3038
timestamp 1681620392
transform 1 0 2212 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3039
timestamp 1681620392
transform 1 0 2276 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3040
timestamp 1681620392
transform 1 0 2308 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3108
timestamp 1681620392
transform 1 0 2196 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3109
timestamp 1681620392
transform 1 0 2228 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2607
timestamp 1681620392
transform 1 0 2268 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_3110
timestamp 1681620392
transform 1 0 2316 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2631
timestamp 1681620392
transform 1 0 2212 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2632
timestamp 1681620392
transform 1 0 2308 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2648
timestamp 1681620392
transform 1 0 2220 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2649
timestamp 1681620392
transform 1 0 2276 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2650
timestamp 1681620392
transform 1 0 2316 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_3111
timestamp 1681620392
transform 1 0 2340 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3112
timestamp 1681620392
transform 1 0 2348 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2633
timestamp 1681620392
transform 1 0 2348 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_3041
timestamp 1681620392
transform 1 0 2396 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_2583
timestamp 1681620392
transform 1 0 2404 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2549
timestamp 1681620392
transform 1 0 2420 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_3042
timestamp 1681620392
transform 1 0 2412 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3113
timestamp 1681620392
transform 1 0 2404 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2651
timestamp 1681620392
transform 1 0 2396 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_3043
timestamp 1681620392
transform 1 0 2436 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3114
timestamp 1681620392
transform 1 0 2428 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2634
timestamp 1681620392
transform 1 0 2428 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2550
timestamp 1681620392
transform 1 0 2460 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_2977
timestamp 1681620392
transform 1 0 2460 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_2584
timestamp 1681620392
transform 1 0 2460 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_3115
timestamp 1681620392
transform 1 0 2452 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3116
timestamp 1681620392
transform 1 0 2460 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2566
timestamp 1681620392
transform 1 0 2492 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2551
timestamp 1681620392
transform 1 0 2516 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_2978
timestamp 1681620392
transform 1 0 2508 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2979
timestamp 1681620392
transform 1 0 2516 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3044
timestamp 1681620392
transform 1 0 2492 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3117
timestamp 1681620392
transform 1 0 2492 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2635
timestamp 1681620392
transform 1 0 2492 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2567
timestamp 1681620392
transform 1 0 2540 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_3045
timestamp 1681620392
transform 1 0 2516 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3046
timestamp 1681620392
transform 1 0 2532 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3047
timestamp 1681620392
transform 1 0 2548 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3118
timestamp 1681620392
transform 1 0 2516 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3119
timestamp 1681620392
transform 1 0 2540 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2585
timestamp 1681620392
transform 1 0 2556 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2533
timestamp 1681620392
transform 1 0 2580 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2568
timestamp 1681620392
transform 1 0 2604 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_3048
timestamp 1681620392
transform 1 0 2580 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3049
timestamp 1681620392
transform 1 0 2588 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_2586
timestamp 1681620392
transform 1 0 2596 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_3050
timestamp 1681620392
transform 1 0 2604 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_2587
timestamp 1681620392
transform 1 0 2612 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_3051
timestamp 1681620392
transform 1 0 2620 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_2588
timestamp 1681620392
transform 1 0 2628 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_3052
timestamp 1681620392
transform 1 0 2668 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_2589
timestamp 1681620392
transform 1 0 2700 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_3120
timestamp 1681620392
transform 1 0 2572 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3121
timestamp 1681620392
transform 1 0 2580 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3122
timestamp 1681620392
transform 1 0 2596 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2608
timestamp 1681620392
transform 1 0 2604 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_3123
timestamp 1681620392
transform 1 0 2612 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2636
timestamp 1681620392
transform 1 0 2588 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2609
timestamp 1681620392
transform 1 0 2652 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2569
timestamp 1681620392
transform 1 0 2732 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2590
timestamp 1681620392
transform 1 0 2724 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2534
timestamp 1681620392
transform 1 0 2756 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_2980
timestamp 1681620392
transform 1 0 2748 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_2570
timestamp 1681620392
transform 1 0 2756 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_3053
timestamp 1681620392
transform 1 0 2732 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3054
timestamp 1681620392
transform 1 0 2740 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3124
timestamp 1681620392
transform 1 0 2700 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3125
timestamp 1681620392
transform 1 0 2716 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3126
timestamp 1681620392
transform 1 0 2732 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2652
timestamp 1681620392
transform 1 0 2700 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_3127
timestamp 1681620392
transform 1 0 2756 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2637
timestamp 1681620392
transform 1 0 2756 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_3128
timestamp 1681620392
transform 1 0 2772 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2638
timestamp 1681620392
transform 1 0 2772 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_3055
timestamp 1681620392
transform 1 0 2780 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3056
timestamp 1681620392
transform 1 0 2788 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_2610
timestamp 1681620392
transform 1 0 2788 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_2981
timestamp 1681620392
transform 1 0 2804 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3057
timestamp 1681620392
transform 1 0 2844 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3129
timestamp 1681620392
transform 1 0 2836 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2653
timestamp 1681620392
transform 1 0 2836 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_3130
timestamp 1681620392
transform 1 0 2868 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3131
timestamp 1681620392
transform 1 0 2876 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_2654
timestamp 1681620392
transform 1 0 2884 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2571
timestamp 1681620392
transform 1 0 2924 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_3058
timestamp 1681620392
transform 1 0 2924 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3132
timestamp 1681620392
transform 1 0 2924 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2982
timestamp 1681620392
transform 1 0 2964 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_2591
timestamp 1681620392
transform 1 0 2956 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2655
timestamp 1681620392
transform 1 0 2972 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_3059
timestamp 1681620392
transform 1 0 3004 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3133
timestamp 1681620392
transform 1 0 2996 0 1 1405
box -2 -2 2 2
use Project_Top_VIA0  Project_Top_VIA0_32
timestamp 1681620392
transform 1 0 48 0 1 1370
box -10 -3 10 3
use FILL  FILL_692
timestamp 1681620392
transform 1 0 72 0 1 1370
box -8 -3 16 105
use FILL  FILL_694
timestamp 1681620392
transform 1 0 80 0 1 1370
box -8 -3 16 105
use FILL  FILL_695
timestamp 1681620392
transform 1 0 88 0 1 1370
box -8 -3 16 105
use FILL  FILL_696
timestamp 1681620392
transform 1 0 96 0 1 1370
box -8 -3 16 105
use FILL  FILL_697
timestamp 1681620392
transform 1 0 104 0 1 1370
box -8 -3 16 105
use FILL  FILL_698
timestamp 1681620392
transform 1 0 112 0 1 1370
box -8 -3 16 105
use FILL  FILL_700
timestamp 1681620392
transform 1 0 120 0 1 1370
box -8 -3 16 105
use FILL  FILL_701
timestamp 1681620392
transform 1 0 128 0 1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_66
timestamp 1681620392
transform 1 0 136 0 1 1370
box -8 -3 32 105
use INVX2  INVX2_198
timestamp 1681620392
transform 1 0 160 0 1 1370
box -9 -3 26 105
use NOR2X1  NOR2X1_67
timestamp 1681620392
transform 1 0 176 0 1 1370
box -8 -3 32 105
use FILL  FILL_702
timestamp 1681620392
transform 1 0 200 0 1 1370
box -8 -3 16 105
use FILL  FILL_703
timestamp 1681620392
transform 1 0 208 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_2656
timestamp 1681620392
transform 1 0 228 0 1 1375
box -3 -3 3 3
use FILL  FILL_704
timestamp 1681620392
transform 1 0 216 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_173
timestamp 1681620392
transform -1 0 248 0 1 1370
box -8 -3 32 105
use FILL  FILL_705
timestamp 1681620392
transform 1 0 248 0 1 1370
box -8 -3 16 105
use FILL  FILL_706
timestamp 1681620392
transform 1 0 256 0 1 1370
box -8 -3 16 105
use FILL  FILL_711
timestamp 1681620392
transform 1 0 264 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_2657
timestamp 1681620392
transform 1 0 284 0 1 1375
box -3 -3 3 3
use NAND2X1  NAND2X1_176
timestamp 1681620392
transform -1 0 296 0 1 1370
box -8 -3 32 105
use M3_M2  M3_M2_2658
timestamp 1681620392
transform 1 0 316 0 1 1375
box -3 -3 3 3
use NAND2X1  NAND2X1_177
timestamp 1681620392
transform -1 0 320 0 1 1370
box -8 -3 32 105
use FILL  FILL_712
timestamp 1681620392
transform 1 0 320 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_178
timestamp 1681620392
transform 1 0 328 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_179
timestamp 1681620392
transform 1 0 352 0 1 1370
box -8 -3 32 105
use FILL  FILL_713
timestamp 1681620392
transform 1 0 376 0 1 1370
box -8 -3 16 105
use FILL  FILL_714
timestamp 1681620392
transform 1 0 384 0 1 1370
box -8 -3 16 105
use FILL  FILL_715
timestamp 1681620392
transform 1 0 392 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_200
timestamp 1681620392
transform -1 0 416 0 1 1370
box -9 -3 26 105
use FILL  FILL_716
timestamp 1681620392
transform 1 0 416 0 1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_64
timestamp 1681620392
transform 1 0 424 0 1 1370
box -8 -3 40 105
use FILL  FILL_717
timestamp 1681620392
transform 1 0 456 0 1 1370
box -8 -3 16 105
use FILL  FILL_718
timestamp 1681620392
transform 1 0 464 0 1 1370
box -8 -3 16 105
use FILL  FILL_719
timestamp 1681620392
transform 1 0 472 0 1 1370
box -8 -3 16 105
use FILL  FILL_720
timestamp 1681620392
transform 1 0 480 0 1 1370
box -8 -3 16 105
use FILL  FILL_721
timestamp 1681620392
transform 1 0 488 0 1 1370
box -8 -3 16 105
use FILL  FILL_722
timestamp 1681620392
transform 1 0 496 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_180
timestamp 1681620392
transform 1 0 504 0 1 1370
box -8 -3 32 105
use FILL  FILL_723
timestamp 1681620392
transform 1 0 528 0 1 1370
box -8 -3 16 105
use FILL  FILL_724
timestamp 1681620392
transform 1 0 536 0 1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_47
timestamp 1681620392
transform -1 0 584 0 1 1370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_177
timestamp 1681620392
transform -1 0 680 0 1 1370
box -8 -3 104 105
use FILL  FILL_725
timestamp 1681620392
transform 1 0 680 0 1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_65
timestamp 1681620392
transform -1 0 720 0 1 1370
box -8 -3 40 105
use INVX2  INVX2_201
timestamp 1681620392
transform 1 0 720 0 1 1370
box -9 -3 26 105
use FILL  FILL_726
timestamp 1681620392
transform 1 0 736 0 1 1370
box -8 -3 16 105
use FILL  FILL_727
timestamp 1681620392
transform 1 0 744 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_181
timestamp 1681620392
transform 1 0 752 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_182
timestamp 1681620392
transform -1 0 800 0 1 1370
box -8 -3 32 105
use FILL  FILL_728
timestamp 1681620392
transform 1 0 800 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_183
timestamp 1681620392
transform 1 0 808 0 1 1370
box -8 -3 32 105
use OAI21X1  OAI21X1_178
timestamp 1681620392
transform 1 0 832 0 1 1370
box -8 -3 34 105
use AND2X2  AND2X2_16
timestamp 1681620392
transform -1 0 896 0 1 1370
box -8 -3 40 105
use FILL  FILL_729
timestamp 1681620392
transform 1 0 896 0 1 1370
box -8 -3 16 105
use FILL  FILL_737
timestamp 1681620392
transform 1 0 904 0 1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_69
timestamp 1681620392
transform 1 0 912 0 1 1370
box -8 -3 40 105
use NAND2X1  NAND2X1_190
timestamp 1681620392
transform -1 0 968 0 1 1370
box -8 -3 32 105
use FILL  FILL_739
timestamp 1681620392
transform 1 0 968 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_180
timestamp 1681620392
transform 1 0 976 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_181
timestamp 1681620392
transform -1 0 1040 0 1 1370
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_179
timestamp 1681620392
transform 1 0 1040 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_207
timestamp 1681620392
transform 1 0 1136 0 1 1370
box -9 -3 26 105
use BUFX2  BUFX2_30
timestamp 1681620392
transform 1 0 1152 0 1 1370
box -5 -3 28 105
use FILL  FILL_744
timestamp 1681620392
transform 1 0 1176 0 1 1370
box -8 -3 16 105
use FILL  FILL_746
timestamp 1681620392
transform 1 0 1184 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_2659
timestamp 1681620392
transform 1 0 1204 0 1 1375
box -3 -3 3 3
use AND2X2  AND2X2_18
timestamp 1681620392
transform 1 0 1192 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_19
timestamp 1681620392
transform 1 0 1224 0 1 1370
box -8 -3 40 105
use FILL  FILL_747
timestamp 1681620392
transform 1 0 1256 0 1 1370
box -8 -3 16 105
use FILL  FILL_750
timestamp 1681620392
transform 1 0 1264 0 1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_70
timestamp 1681620392
transform 1 0 1272 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_71
timestamp 1681620392
transform 1 0 1304 0 1 1370
box -8 -3 40 105
use M3_M2  M3_M2_2660
timestamp 1681620392
transform 1 0 1364 0 1 1375
box -3 -3 3 3
use INVX2  INVX2_209
timestamp 1681620392
transform 1 0 1336 0 1 1370
box -9 -3 26 105
use OAI21X1  OAI21X1_185
timestamp 1681620392
transform 1 0 1352 0 1 1370
box -8 -3 34 105
use FILL  FILL_751
timestamp 1681620392
transform 1 0 1384 0 1 1370
box -8 -3 16 105
use FILL  FILL_752
timestamp 1681620392
transform 1 0 1392 0 1 1370
box -8 -3 16 105
use FILL  FILL_759
timestamp 1681620392
transform 1 0 1400 0 1 1370
box -8 -3 16 105
use FILL  FILL_761
timestamp 1681620392
transform 1 0 1408 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_192
timestamp 1681620392
transform -1 0 1440 0 1 1370
box -8 -3 32 105
use FILL  FILL_762
timestamp 1681620392
transform 1 0 1440 0 1 1370
box -8 -3 16 105
use FILL  FILL_763
timestamp 1681620392
transform 1 0 1448 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_193
timestamp 1681620392
transform 1 0 1456 0 1 1370
box -8 -3 32 105
use OAI22X1  OAI22X1_50
timestamp 1681620392
transform -1 0 1520 0 1 1370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_181
timestamp 1681620392
transform -1 0 1616 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_182
timestamp 1681620392
transform -1 0 1712 0 1 1370
box -8 -3 104 105
use BUFX2  BUFX2_33
timestamp 1681620392
transform 1 0 1712 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_34
timestamp 1681620392
transform 1 0 1736 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_35
timestamp 1681620392
transform 1 0 1760 0 1 1370
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_183
timestamp 1681620392
transform 1 0 1784 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_210
timestamp 1681620392
transform 1 0 1880 0 1 1370
box -9 -3 26 105
use FILL  FILL_764
timestamp 1681620392
transform 1 0 1896 0 1 1370
box -8 -3 16 105
use FILL  FILL_765
timestamp 1681620392
transform 1 0 1904 0 1 1370
box -8 -3 16 105
use FILL  FILL_766
timestamp 1681620392
transform 1 0 1912 0 1 1370
box -8 -3 16 105
use FILL  FILL_767
timestamp 1681620392
transform 1 0 1920 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_186
timestamp 1681620392
transform 1 0 1928 0 1 1370
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_184
timestamp 1681620392
transform 1 0 1960 0 1 1370
box -8 -3 104 105
use FILL  FILL_768
timestamp 1681620392
transform 1 0 2056 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_194
timestamp 1681620392
transform 1 0 2064 0 1 1370
box -8 -3 32 105
use INVX2  INVX2_211
timestamp 1681620392
transform 1 0 2088 0 1 1370
box -9 -3 26 105
use NAND2X1  NAND2X1_195
timestamp 1681620392
transform 1 0 2104 0 1 1370
box -8 -3 32 105
use M3_M2  M3_M2_2661
timestamp 1681620392
transform 1 0 2140 0 1 1375
box -3 -3 3 3
use FILL  FILL_769
timestamp 1681620392
transform 1 0 2128 0 1 1370
box -8 -3 16 105
use FILL  FILL_770
timestamp 1681620392
transform 1 0 2136 0 1 1370
box -8 -3 16 105
use FILL  FILL_771
timestamp 1681620392
transform 1 0 2144 0 1 1370
box -8 -3 16 105
use FILL  FILL_772
timestamp 1681620392
transform 1 0 2152 0 1 1370
box -8 -3 16 105
use FILL  FILL_773
timestamp 1681620392
transform 1 0 2160 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_187
timestamp 1681620392
transform 1 0 2168 0 1 1370
box -8 -3 34 105
use INVX2  INVX2_212
timestamp 1681620392
transform 1 0 2200 0 1 1370
box -9 -3 26 105
use M3_M2  M3_M2_2662
timestamp 1681620392
transform 1 0 2284 0 1 1375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_185
timestamp 1681620392
transform 1 0 2216 0 1 1370
box -8 -3 104 105
use M3_M2  M3_M2_2663
timestamp 1681620392
transform 1 0 2332 0 1 1375
box -3 -3 3 3
use OAI21X1  OAI21X1_188
timestamp 1681620392
transform -1 0 2344 0 1 1370
box -8 -3 34 105
use INVX2  INVX2_213
timestamp 1681620392
transform 1 0 2344 0 1 1370
box -9 -3 26 105
use FILL  FILL_774
timestamp 1681620392
transform 1 0 2360 0 1 1370
box -8 -3 16 105
use FILL  FILL_775
timestamp 1681620392
transform 1 0 2368 0 1 1370
box -8 -3 16 105
use FILL  FILL_776
timestamp 1681620392
transform 1 0 2376 0 1 1370
box -8 -3 16 105
use FILL  FILL_777
timestamp 1681620392
transform 1 0 2384 0 1 1370
box -8 -3 16 105
use FILL  FILL_778
timestamp 1681620392
transform 1 0 2392 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_2664
timestamp 1681620392
transform 1 0 2428 0 1 1375
box -3 -3 3 3
use NAND2X1  NAND2X1_196
timestamp 1681620392
transform 1 0 2400 0 1 1370
box -8 -3 32 105
use OAI21X1  OAI21X1_189
timestamp 1681620392
transform 1 0 2424 0 1 1370
box -8 -3 34 105
use FILL  FILL_779
timestamp 1681620392
transform 1 0 2456 0 1 1370
box -8 -3 16 105
use FILL  FILL_780
timestamp 1681620392
transform 1 0 2464 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_214
timestamp 1681620392
transform 1 0 2472 0 1 1370
box -9 -3 26 105
use M3_M2  M3_M2_2665
timestamp 1681620392
transform 1 0 2524 0 1 1375
box -3 -3 3 3
use NAND2X1  NAND2X1_197
timestamp 1681620392
transform 1 0 2488 0 1 1370
box -8 -3 32 105
use OAI21X1  OAI21X1_190
timestamp 1681620392
transform -1 0 2544 0 1 1370
box -8 -3 34 105
use FILL  FILL_781
timestamp 1681620392
transform 1 0 2544 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_2666
timestamp 1681620392
transform 1 0 2580 0 1 1375
box -3 -3 3 3
use BUFX2  BUFX2_36
timestamp 1681620392
transform 1 0 2552 0 1 1370
box -5 -3 28 105
use OAI22X1  OAI22X1_51
timestamp 1681620392
transform 1 0 2576 0 1 1370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_186
timestamp 1681620392
transform -1 0 2712 0 1 1370
box -8 -3 104 105
use M3_M2  M3_M2_2667
timestamp 1681620392
transform 1 0 2724 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2668
timestamp 1681620392
transform 1 0 2740 0 1 1375
box -3 -3 3 3
use INVX2  INVX2_215
timestamp 1681620392
transform 1 0 2712 0 1 1370
box -9 -3 26 105
use NAND2X1  NAND2X1_198
timestamp 1681620392
transform 1 0 2728 0 1 1370
box -8 -3 32 105
use M3_M2  M3_M2_2669
timestamp 1681620392
transform 1 0 2772 0 1 1375
box -3 -3 3 3
use INVX2  INVX2_222
timestamp 1681620392
transform 1 0 2752 0 1 1370
box -9 -3 26 105
use FILL  FILL_785
timestamp 1681620392
transform 1 0 2768 0 1 1370
box -8 -3 16 105
use FILL  FILL_786
timestamp 1681620392
transform 1 0 2776 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_204
timestamp 1681620392
transform 1 0 2784 0 1 1370
box -8 -3 32 105
use FILL  FILL_787
timestamp 1681620392
transform 1 0 2808 0 1 1370
box -8 -3 16 105
use FILL  FILL_789
timestamp 1681620392
transform 1 0 2816 0 1 1370
box -8 -3 16 105
use FILL  FILL_791
timestamp 1681620392
transform 1 0 2824 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_198
timestamp 1681620392
transform 1 0 2832 0 1 1370
box -8 -3 34 105
use FILL  FILL_793
timestamp 1681620392
transform 1 0 2864 0 1 1370
box -8 -3 16 105
use FILL  FILL_794
timestamp 1681620392
transform 1 0 2872 0 1 1370
box -8 -3 16 105
use FILL  FILL_796
timestamp 1681620392
transform 1 0 2880 0 1 1370
box -8 -3 16 105
use FILL  FILL_798
timestamp 1681620392
transform 1 0 2888 0 1 1370
box -8 -3 16 105
use FILL  FILL_800
timestamp 1681620392
transform 1 0 2896 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_223
timestamp 1681620392
transform 1 0 2904 0 1 1370
box -9 -3 26 105
use NAND2X1  NAND2X1_206
timestamp 1681620392
transform 1 0 2920 0 1 1370
box -8 -3 32 105
use FILL  FILL_802
timestamp 1681620392
transform 1 0 2944 0 1 1370
box -8 -3 16 105
use FILL  FILL_804
timestamp 1681620392
transform 1 0 2952 0 1 1370
box -8 -3 16 105
use FILL  FILL_806
timestamp 1681620392
transform 1 0 2960 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_199
timestamp 1681620392
transform -1 0 3000 0 1 1370
box -8 -3 34 105
use FILL  FILL_807
timestamp 1681620392
transform 1 0 3000 0 1 1370
box -8 -3 16 105
use FILL  FILL_812
timestamp 1681620392
transform 1 0 3008 0 1 1370
box -8 -3 16 105
use Project_Top_VIA0  Project_Top_VIA0_33
timestamp 1681620392
transform 1 0 3043 0 1 1370
box -10 -3 10 3
use M2_M1  M2_M1_3141
timestamp 1681620392
transform 1 0 92 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3224
timestamp 1681620392
transform 1 0 84 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2757
timestamp 1681620392
transform 1 0 92 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_3225
timestamp 1681620392
transform 1 0 108 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2780
timestamp 1681620392
transform 1 0 84 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2670
timestamp 1681620392
transform 1 0 140 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2691
timestamp 1681620392
transform 1 0 164 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2692
timestamp 1681620392
transform 1 0 180 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_3136
timestamp 1681620392
transform 1 0 148 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_2714
timestamp 1681620392
transform 1 0 156 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3137
timestamp 1681620392
transform 1 0 188 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_3142
timestamp 1681620392
transform 1 0 140 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3143
timestamp 1681620392
transform 1 0 156 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3144
timestamp 1681620392
transform 1 0 172 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3145
timestamp 1681620392
transform 1 0 180 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3226
timestamp 1681620392
transform 1 0 172 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2671
timestamp 1681620392
transform 1 0 204 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_3227
timestamp 1681620392
transform 1 0 188 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2830
timestamp 1681620392
transform 1 0 180 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2758
timestamp 1681620392
transform 1 0 196 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_3310
timestamp 1681620392
transform 1 0 196 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2742
timestamp 1681620392
transform 1 0 212 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_3146
timestamp 1681620392
transform 1 0 228 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3147
timestamp 1681620392
transform 1 0 236 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_2715
timestamp 1681620392
transform 1 0 252 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3148
timestamp 1681620392
transform 1 0 252 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_2743
timestamp 1681620392
transform 1 0 260 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_3228
timestamp 1681620392
transform 1 0 244 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2781
timestamp 1681620392
transform 1 0 236 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2759
timestamp 1681620392
transform 1 0 252 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_3229
timestamp 1681620392
transform 1 0 260 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3311
timestamp 1681620392
transform 1 0 252 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2810
timestamp 1681620392
transform 1 0 252 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2811
timestamp 1681620392
transform 1 0 268 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2852
timestamp 1681620392
transform 1 0 276 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_3312
timestamp 1681620392
transform 1 0 292 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3313
timestamp 1681620392
transform 1 0 300 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2831
timestamp 1681620392
transform 1 0 300 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2853
timestamp 1681620392
transform 1 0 292 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_3138
timestamp 1681620392
transform 1 0 356 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_3149
timestamp 1681620392
transform 1 0 340 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3230
timestamp 1681620392
transform 1 0 316 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3231
timestamp 1681620392
transform 1 0 324 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3232
timestamp 1681620392
transform 1 0 356 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3233
timestamp 1681620392
transform 1 0 364 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2782
timestamp 1681620392
transform 1 0 324 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2783
timestamp 1681620392
transform 1 0 340 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2832
timestamp 1681620392
transform 1 0 316 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2716
timestamp 1681620392
transform 1 0 388 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3139
timestamp 1681620392
transform 1 0 404 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_3150
timestamp 1681620392
transform 1 0 372 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3151
timestamp 1681620392
transform 1 0 388 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3234
timestamp 1681620392
transform 1 0 372 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3235
timestamp 1681620392
transform 1 0 380 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2784
timestamp 1681620392
transform 1 0 372 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_3152
timestamp 1681620392
transform 1 0 444 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3153
timestamp 1681620392
transform 1 0 460 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3236
timestamp 1681620392
transform 1 0 404 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2760
timestamp 1681620392
transform 1 0 412 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_3237
timestamp 1681620392
transform 1 0 420 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2761
timestamp 1681620392
transform 1 0 428 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_3238
timestamp 1681620392
transform 1 0 444 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3314
timestamp 1681620392
transform 1 0 412 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2812
timestamp 1681620392
transform 1 0 404 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_3343
timestamp 1681620392
transform 1 0 412 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_3315
timestamp 1681620392
transform 1 0 436 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2833
timestamp 1681620392
transform 1 0 420 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_3239
timestamp 1681620392
transform 1 0 468 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2762
timestamp 1681620392
transform 1 0 476 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_3316
timestamp 1681620392
transform 1 0 476 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3317
timestamp 1681620392
transform 1 0 484 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2813
timestamp 1681620392
transform 1 0 484 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2834
timestamp 1681620392
transform 1 0 468 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_3154
timestamp 1681620392
transform 1 0 500 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3240
timestamp 1681620392
transform 1 0 500 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2763
timestamp 1681620392
transform 1 0 508 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2785
timestamp 1681620392
transform 1 0 500 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_3318
timestamp 1681620392
transform 1 0 508 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3155
timestamp 1681620392
transform 1 0 524 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_2764
timestamp 1681620392
transform 1 0 532 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2693
timestamp 1681620392
transform 1 0 588 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_3156
timestamp 1681620392
transform 1 0 556 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_2744
timestamp 1681620392
transform 1 0 564 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2717
timestamp 1681620392
transform 1 0 604 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2718
timestamp 1681620392
transform 1 0 652 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3157
timestamp 1681620392
transform 1 0 588 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3158
timestamp 1681620392
transform 1 0 604 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3241
timestamp 1681620392
transform 1 0 540 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3242
timestamp 1681620392
transform 1 0 564 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3243
timestamp 1681620392
transform 1 0 580 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2786
timestamp 1681620392
transform 1 0 540 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2787
timestamp 1681620392
transform 1 0 564 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2835
timestamp 1681620392
transform 1 0 556 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2745
timestamp 1681620392
transform 1 0 628 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2765
timestamp 1681620392
transform 1 0 604 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_3244
timestamp 1681620392
transform 1 0 628 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2766
timestamp 1681620392
transform 1 0 636 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2854
timestamp 1681620392
transform 1 0 596 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_3159
timestamp 1681620392
transform 1 0 708 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3160
timestamp 1681620392
transform 1 0 724 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3161
timestamp 1681620392
transform 1 0 740 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3162
timestamp 1681620392
transform 1 0 756 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3163
timestamp 1681620392
transform 1 0 772 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3245
timestamp 1681620392
transform 1 0 700 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3246
timestamp 1681620392
transform 1 0 716 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3247
timestamp 1681620392
transform 1 0 732 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3248
timestamp 1681620392
transform 1 0 748 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2788
timestamp 1681620392
transform 1 0 716 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2789
timestamp 1681620392
transform 1 0 748 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_3319
timestamp 1681620392
transform 1 0 764 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3249
timestamp 1681620392
transform 1 0 796 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3320
timestamp 1681620392
transform 1 0 788 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3344
timestamp 1681620392
transform 1 0 780 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_3250
timestamp 1681620392
transform 1 0 828 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3348
timestamp 1681620392
transform 1 0 828 0 1 1295
box -2 -2 2 2
use M2_M1  M2_M1_3164
timestamp 1681620392
transform 1 0 852 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_2746
timestamp 1681620392
transform 1 0 860 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_3321
timestamp 1681620392
transform 1 0 860 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3345
timestamp 1681620392
transform 1 0 844 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_2814
timestamp 1681620392
transform 1 0 860 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2694
timestamp 1681620392
transform 1 0 892 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_3165
timestamp 1681620392
transform 1 0 884 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3322
timestamp 1681620392
transform 1 0 884 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2747
timestamp 1681620392
transform 1 0 900 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2815
timestamp 1681620392
transform 1 0 900 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_3251
timestamp 1681620392
transform 1 0 924 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2790
timestamp 1681620392
transform 1 0 924 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_3166
timestamp 1681620392
transform 1 0 940 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3252
timestamp 1681620392
transform 1 0 948 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2695
timestamp 1681620392
transform 1 0 996 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_3167
timestamp 1681620392
transform 1 0 972 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3168
timestamp 1681620392
transform 1 0 988 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3169
timestamp 1681620392
transform 1 0 996 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3253
timestamp 1681620392
transform 1 0 964 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3254
timestamp 1681620392
transform 1 0 980 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2791
timestamp 1681620392
transform 1 0 964 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2672
timestamp 1681620392
transform 1 0 1052 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2673
timestamp 1681620392
transform 1 0 1092 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2696
timestamp 1681620392
transform 1 0 1036 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2719
timestamp 1681620392
transform 1 0 1028 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2720
timestamp 1681620392
transform 1 0 1068 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2748
timestamp 1681620392
transform 1 0 1012 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_3170
timestamp 1681620392
transform 1 0 1028 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3171
timestamp 1681620392
transform 1 0 1044 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3255
timestamp 1681620392
transform 1 0 1012 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2749
timestamp 1681620392
transform 1 0 1076 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_3172
timestamp 1681620392
transform 1 0 1132 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3256
timestamp 1681620392
transform 1 0 1068 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3257
timestamp 1681620392
transform 1 0 1124 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3258
timestamp 1681620392
transform 1 0 1148 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3323
timestamp 1681620392
transform 1 0 1028 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2836
timestamp 1681620392
transform 1 0 1012 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2837
timestamp 1681620392
transform 1 0 1044 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2838
timestamp 1681620392
transform 1 0 1116 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2674
timestamp 1681620392
transform 1 0 1172 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2697
timestamp 1681620392
transform 1 0 1172 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_3173
timestamp 1681620392
transform 1 0 1172 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_2675
timestamp 1681620392
transform 1 0 1204 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_3174
timestamp 1681620392
transform 1 0 1212 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3259
timestamp 1681620392
transform 1 0 1196 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3324
timestamp 1681620392
transform 1 0 1228 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2816
timestamp 1681620392
transform 1 0 1228 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_3175
timestamp 1681620392
transform 1 0 1268 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3325
timestamp 1681620392
transform 1 0 1276 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3176
timestamp 1681620392
transform 1 0 1300 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_2767
timestamp 1681620392
transform 1 0 1292 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_3326
timestamp 1681620392
transform 1 0 1292 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3346
timestamp 1681620392
transform 1 0 1300 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_3260
timestamp 1681620392
transform 1 0 1324 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2792
timestamp 1681620392
transform 1 0 1324 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2721
timestamp 1681620392
transform 1 0 1364 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3327
timestamp 1681620392
transform 1 0 1348 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2793
timestamp 1681620392
transform 1 0 1356 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_3261
timestamp 1681620392
transform 1 0 1372 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3328
timestamp 1681620392
transform 1 0 1364 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3329
timestamp 1681620392
transform 1 0 1388 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3347
timestamp 1681620392
transform 1 0 1380 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_2722
timestamp 1681620392
transform 1 0 1412 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3177
timestamp 1681620392
transform 1 0 1404 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_2768
timestamp 1681620392
transform 1 0 1420 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2769
timestamp 1681620392
transform 1 0 1444 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2698
timestamp 1681620392
transform 1 0 1500 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2699
timestamp 1681620392
transform 1 0 1516 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2723
timestamp 1681620392
transform 1 0 1492 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3178
timestamp 1681620392
transform 1 0 1484 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3179
timestamp 1681620392
transform 1 0 1492 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3262
timestamp 1681620392
transform 1 0 1460 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3263
timestamp 1681620392
transform 1 0 1476 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3330
timestamp 1681620392
transform 1 0 1444 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2817
timestamp 1681620392
transform 1 0 1436 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2855
timestamp 1681620392
transform 1 0 1428 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2770
timestamp 1681620392
transform 1 0 1484 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_3264
timestamp 1681620392
transform 1 0 1492 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3331
timestamp 1681620392
transform 1 0 1476 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2818
timestamp 1681620392
transform 1 0 1476 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2839
timestamp 1681620392
transform 1 0 1460 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2794
timestamp 1681620392
transform 1 0 1492 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2724
timestamp 1681620392
transform 1 0 1516 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3180
timestamp 1681620392
transform 1 0 1516 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_2771
timestamp 1681620392
transform 1 0 1516 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2676
timestamp 1681620392
transform 1 0 1548 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2677
timestamp 1681620392
transform 1 0 1604 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2700
timestamp 1681620392
transform 1 0 1564 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2701
timestamp 1681620392
transform 1 0 1588 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2725
timestamp 1681620392
transform 1 0 1572 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3181
timestamp 1681620392
transform 1 0 1532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3182
timestamp 1681620392
transform 1 0 1548 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3265
timestamp 1681620392
transform 1 0 1524 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3332
timestamp 1681620392
transform 1 0 1516 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2840
timestamp 1681620392
transform 1 0 1508 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2841
timestamp 1681620392
transform 1 0 1524 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_3266
timestamp 1681620392
transform 1 0 1572 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2856
timestamp 1681620392
transform 1 0 1548 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_3183
timestamp 1681620392
transform 1 0 1652 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3267
timestamp 1681620392
transform 1 0 1644 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2795
timestamp 1681620392
transform 1 0 1644 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2726
timestamp 1681620392
transform 1 0 1668 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3184
timestamp 1681620392
transform 1 0 1668 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3185
timestamp 1681620392
transform 1 0 1692 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_2772
timestamp 1681620392
transform 1 0 1684 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_3333
timestamp 1681620392
transform 1 0 1692 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2678
timestamp 1681620392
transform 1 0 1732 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2702
timestamp 1681620392
transform 1 0 1716 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2703
timestamp 1681620392
transform 1 0 1756 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2727
timestamp 1681620392
transform 1 0 1716 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3186
timestamp 1681620392
transform 1 0 1716 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3187
timestamp 1681620392
transform 1 0 1732 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3268
timestamp 1681620392
transform 1 0 1716 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3269
timestamp 1681620392
transform 1 0 1780 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2796
timestamp 1681620392
transform 1 0 1780 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2819
timestamp 1681620392
transform 1 0 1716 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2679
timestamp 1681620392
transform 1 0 1940 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2680
timestamp 1681620392
transform 1 0 1964 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2728
timestamp 1681620392
transform 1 0 1884 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3188
timestamp 1681620392
transform 1 0 1836 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3189
timestamp 1681620392
transform 1 0 1852 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3190
timestamp 1681620392
transform 1 0 1868 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3191
timestamp 1681620392
transform 1 0 1884 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3270
timestamp 1681620392
transform 1 0 1828 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3271
timestamp 1681620392
transform 1 0 1844 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2773
timestamp 1681620392
transform 1 0 1852 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_3272
timestamp 1681620392
transform 1 0 1860 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2797
timestamp 1681620392
transform 1 0 1844 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2820
timestamp 1681620392
transform 1 0 1860 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2774
timestamp 1681620392
transform 1 0 1916 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2704
timestamp 1681620392
transform 1 0 2020 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2705
timestamp 1681620392
transform 1 0 2068 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2729
timestamp 1681620392
transform 1 0 2004 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2730
timestamp 1681620392
transform 1 0 2052 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3192
timestamp 1681620392
transform 1 0 1988 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3193
timestamp 1681620392
transform 1 0 2004 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3273
timestamp 1681620392
transform 1 0 1924 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3274
timestamp 1681620392
transform 1 0 1972 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3275
timestamp 1681620392
transform 1 0 1980 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2798
timestamp 1681620392
transform 1 0 1932 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_3334
timestamp 1681620392
transform 1 0 1972 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2799
timestamp 1681620392
transform 1 0 1980 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2821
timestamp 1681620392
transform 1 0 1980 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2731
timestamp 1681620392
transform 1 0 2108 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2681
timestamp 1681620392
transform 1 0 2140 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_3194
timestamp 1681620392
transform 1 0 2108 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3195
timestamp 1681620392
transform 1 0 2124 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3196
timestamp 1681620392
transform 1 0 2148 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3276
timestamp 1681620392
transform 1 0 2052 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3277
timestamp 1681620392
transform 1 0 2084 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3278
timestamp 1681620392
transform 1 0 2092 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3279
timestamp 1681620392
transform 1 0 2100 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3280
timestamp 1681620392
transform 1 0 2116 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2775
timestamp 1681620392
transform 1 0 2124 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2706
timestamp 1681620392
transform 1 0 2228 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_3197
timestamp 1681620392
transform 1 0 2180 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3281
timestamp 1681620392
transform 1 0 2140 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3282
timestamp 1681620392
transform 1 0 2156 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3283
timestamp 1681620392
transform 1 0 2164 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3284
timestamp 1681620392
transform 1 0 2204 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3285
timestamp 1681620392
transform 1 0 2260 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3286
timestamp 1681620392
transform 1 0 2276 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2800
timestamp 1681620392
transform 1 0 2044 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2801
timestamp 1681620392
transform 1 0 2084 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2822
timestamp 1681620392
transform 1 0 2092 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2842
timestamp 1681620392
transform 1 0 2004 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2843
timestamp 1681620392
transform 1 0 2044 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2823
timestamp 1681620392
transform 1 0 2164 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2844
timestamp 1681620392
transform 1 0 2252 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2682
timestamp 1681620392
transform 1 0 2356 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2707
timestamp 1681620392
transform 1 0 2300 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_3198
timestamp 1681620392
transform 1 0 2300 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_2750
timestamp 1681620392
transform 1 0 2340 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_3287
timestamp 1681620392
transform 1 0 2324 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3335
timestamp 1681620392
transform 1 0 2284 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2824
timestamp 1681620392
transform 1 0 2276 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2845
timestamp 1681620392
transform 1 0 2276 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2857
timestamp 1681620392
transform 1 0 2284 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2858
timestamp 1681620392
transform 1 0 2316 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2708
timestamp 1681620392
transform 1 0 2404 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2732
timestamp 1681620392
transform 1 0 2436 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3199
timestamp 1681620392
transform 1 0 2404 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3200
timestamp 1681620392
transform 1 0 2428 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3288
timestamp 1681620392
transform 1 0 2396 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3289
timestamp 1681620392
transform 1 0 2412 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3336
timestamp 1681620392
transform 1 0 2428 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3201
timestamp 1681620392
transform 1 0 2436 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_2751
timestamp 1681620392
transform 1 0 2452 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2683
timestamp 1681620392
transform 1 0 2492 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2684
timestamp 1681620392
transform 1 0 2516 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2685
timestamp 1681620392
transform 1 0 2540 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_3202
timestamp 1681620392
transform 1 0 2468 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_2709
timestamp 1681620392
transform 1 0 2508 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2733
timestamp 1681620392
transform 1 0 2516 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2734
timestamp 1681620392
transform 1 0 2564 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2686
timestamp 1681620392
transform 1 0 2612 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2735
timestamp 1681620392
transform 1 0 2588 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3203
timestamp 1681620392
transform 1 0 2492 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3204
timestamp 1681620392
transform 1 0 2580 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3205
timestamp 1681620392
transform 1 0 2596 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_2752
timestamp 1681620392
transform 1 0 2604 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2710
timestamp 1681620392
transform 1 0 2628 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_3206
timestamp 1681620392
transform 1 0 2612 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3207
timestamp 1681620392
transform 1 0 2620 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3290
timestamp 1681620392
transform 1 0 2452 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3291
timestamp 1681620392
transform 1 0 2460 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3292
timestamp 1681620392
transform 1 0 2476 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3293
timestamp 1681620392
transform 1 0 2516 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3294
timestamp 1681620392
transform 1 0 2572 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3295
timestamp 1681620392
transform 1 0 2588 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3296
timestamp 1681620392
transform 1 0 2604 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3337
timestamp 1681620392
transform 1 0 2436 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2802
timestamp 1681620392
transform 1 0 2460 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2825
timestamp 1681620392
transform 1 0 2436 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2826
timestamp 1681620392
transform 1 0 2476 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2803
timestamp 1681620392
transform 1 0 2604 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2753
timestamp 1681620392
transform 1 0 2636 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2687
timestamp 1681620392
transform 1 0 2692 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2711
timestamp 1681620392
transform 1 0 2660 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2712
timestamp 1681620392
transform 1 0 2716 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2736
timestamp 1681620392
transform 1 0 2684 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2737
timestamp 1681620392
transform 1 0 2708 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3208
timestamp 1681620392
transform 1 0 2652 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3209
timestamp 1681620392
transform 1 0 2668 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_2754
timestamp 1681620392
transform 1 0 2676 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_3210
timestamp 1681620392
transform 1 0 2684 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3211
timestamp 1681620392
transform 1 0 2692 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3212
timestamp 1681620392
transform 1 0 2708 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3297
timestamp 1681620392
transform 1 0 2636 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3298
timestamp 1681620392
transform 1 0 2644 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2776
timestamp 1681620392
transform 1 0 2652 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2755
timestamp 1681620392
transform 1 0 2716 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2688
timestamp 1681620392
transform 1 0 2740 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_3213
timestamp 1681620392
transform 1 0 2724 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3214
timestamp 1681620392
transform 1 0 2732 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3299
timestamp 1681620392
transform 1 0 2660 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3300
timestamp 1681620392
transform 1 0 2676 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3338
timestamp 1681620392
transform 1 0 2620 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2804
timestamp 1681620392
transform 1 0 2628 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2846
timestamp 1681620392
transform 1 0 2620 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2777
timestamp 1681620392
transform 1 0 2692 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2738
timestamp 1681620392
transform 1 0 2748 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3215
timestamp 1681620392
transform 1 0 2756 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3301
timestamp 1681620392
transform 1 0 2700 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3302
timestamp 1681620392
transform 1 0 2716 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2805
timestamp 1681620392
transform 1 0 2676 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2778
timestamp 1681620392
transform 1 0 2732 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_3303
timestamp 1681620392
transform 1 0 2740 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3304
timestamp 1681620392
transform 1 0 2748 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2827
timestamp 1681620392
transform 1 0 2716 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2847
timestamp 1681620392
transform 1 0 2668 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2848
timestamp 1681620392
transform 1 0 2684 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2713
timestamp 1681620392
transform 1 0 2804 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_3216
timestamp 1681620392
transform 1 0 2780 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3217
timestamp 1681620392
transform 1 0 2788 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3339
timestamp 1681620392
transform 1 0 2748 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2806
timestamp 1681620392
transform 1 0 2772 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_3340
timestamp 1681620392
transform 1 0 2780 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2828
timestamp 1681620392
transform 1 0 2748 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_3218
timestamp 1681620392
transform 1 0 2812 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3341
timestamp 1681620392
transform 1 0 2804 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2829
timestamp 1681620392
transform 1 0 2788 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2849
timestamp 1681620392
transform 1 0 2780 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2779
timestamp 1681620392
transform 1 0 2820 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_3342
timestamp 1681620392
transform 1 0 2820 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_2850
timestamp 1681620392
transform 1 0 2812 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2689
timestamp 1681620392
transform 1 0 2836 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2739
timestamp 1681620392
transform 1 0 2852 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2690
timestamp 1681620392
transform 1 0 2876 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_3140
timestamp 1681620392
transform 1 0 2876 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_3219
timestamp 1681620392
transform 1 0 2836 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3220
timestamp 1681620392
transform 1 0 2852 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3221
timestamp 1681620392
transform 1 0 2868 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3305
timestamp 1681620392
transform 1 0 2836 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3306
timestamp 1681620392
transform 1 0 2860 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2807
timestamp 1681620392
transform 1 0 2852 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2756
timestamp 1681620392
transform 1 0 2876 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_3222
timestamp 1681620392
transform 1 0 2916 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_2808
timestamp 1681620392
transform 1 0 2908 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2740
timestamp 1681620392
transform 1 0 2940 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3307
timestamp 1681620392
transform 1 0 2924 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3308
timestamp 1681620392
transform 1 0 2932 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_2809
timestamp 1681620392
transform 1 0 2932 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2851
timestamp 1681620392
transform 1 0 2924 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_3223
timestamp 1681620392
transform 1 0 2948 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_2741
timestamp 1681620392
transform 1 0 2996 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_3309
timestamp 1681620392
transform 1 0 3004 0 1 1325
box -2 -2 2 2
use Project_Top_VIA0  Project_Top_VIA0_34
timestamp 1681620392
transform 1 0 24 0 1 1270
box -10 -3 10 3
use FILL  FILL_693
timestamp 1681620392
transform 1 0 72 0 -1 1370
box -8 -3 16 105
use AOI21X1  AOI21X1_18
timestamp 1681620392
transform 1 0 80 0 -1 1370
box -7 -3 39 105
use FILL  FILL_699
timestamp 1681620392
transform 1 0 112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_707
timestamp 1681620392
transform 1 0 120 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_199
timestamp 1681620392
transform -1 0 144 0 -1 1370
box -9 -3 26 105
use NOR2X1  NOR2X1_68
timestamp 1681620392
transform 1 0 144 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_69
timestamp 1681620392
transform -1 0 192 0 -1 1370
box -8 -3 32 105
use FILL  FILL_708
timestamp 1681620392
transform 1 0 192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_709
timestamp 1681620392
transform 1 0 200 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_2859
timestamp 1681620392
transform 1 0 236 0 1 1275
box -3 -3 3 3
use NAND2X1  NAND2X1_174
timestamp 1681620392
transform -1 0 232 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_175
timestamp 1681620392
transform 1 0 232 0 -1 1370
box -8 -3 32 105
use FILL  FILL_710
timestamp 1681620392
transform 1 0 256 0 -1 1370
box -8 -3 16 105
use FILL  FILL_730
timestamp 1681620392
transform 1 0 264 0 -1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_184
timestamp 1681620392
transform 1 0 272 0 -1 1370
box -8 -3 32 105
use M3_M2  M3_M2_2860
timestamp 1681620392
transform 1 0 308 0 1 1275
box -3 -3 3 3
use FILL  FILL_731
timestamp 1681620392
transform 1 0 296 0 -1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_185
timestamp 1681620392
transform -1 0 328 0 -1 1370
box -8 -3 32 105
use AOI21X1  AOI21X1_19
timestamp 1681620392
transform 1 0 328 0 -1 1370
box -7 -3 39 105
use INVX2  INVX2_202
timestamp 1681620392
transform -1 0 376 0 -1 1370
box -9 -3 26 105
use AOI21X1  AOI21X1_20
timestamp 1681620392
transform 1 0 376 0 -1 1370
box -7 -3 39 105
use NAND3X1  NAND3X1_66
timestamp 1681620392
transform 1 0 408 0 -1 1370
box -8 -3 40 105
use INVX2  INVX2_203
timestamp 1681620392
transform 1 0 440 0 -1 1370
box -9 -3 26 105
use NAND2X1  NAND2X1_186
timestamp 1681620392
transform 1 0 456 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_187
timestamp 1681620392
transform -1 0 504 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_188
timestamp 1681620392
transform -1 0 528 0 -1 1370
box -8 -3 32 105
use OAI21X1  OAI21X1_179
timestamp 1681620392
transform 1 0 528 0 -1 1370
box -8 -3 34 105
use M3_M2  M3_M2_2861
timestamp 1681620392
transform 1 0 580 0 1 1275
box -3 -3 3 3
use AND2X2  AND2X2_17
timestamp 1681620392
transform -1 0 592 0 -1 1370
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_178
timestamp 1681620392
transform 1 0 592 0 -1 1370
box -8 -3 104 105
use INVX2  INVX2_204
timestamp 1681620392
transform 1 0 688 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_205
timestamp 1681620392
transform 1 0 704 0 -1 1370
box -9 -3 26 105
use OAI22X1  OAI22X1_48
timestamp 1681620392
transform -1 0 760 0 -1 1370
box -8 -3 46 105
use NAND3X1  NAND3X1_67
timestamp 1681620392
transform 1 0 760 0 -1 1370
box -8 -3 40 105
use INVX2  INVX2_206
timestamp 1681620392
transform 1 0 792 0 -1 1370
box -9 -3 26 105
use FILL  FILL_732
timestamp 1681620392
transform 1 0 808 0 -1 1370
box -8 -3 16 105
use FILL  FILL_733
timestamp 1681620392
transform 1 0 816 0 -1 1370
box -8 -3 16 105
use FILL  FILL_734
timestamp 1681620392
transform 1 0 824 0 -1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_68
timestamp 1681620392
transform -1 0 864 0 -1 1370
box -8 -3 40 105
use NAND2X1  NAND2X1_189
timestamp 1681620392
transform 1 0 864 0 -1 1370
box -8 -3 32 105
use FILL  FILL_735
timestamp 1681620392
transform 1 0 888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_736
timestamp 1681620392
transform 1 0 896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_738
timestamp 1681620392
transform 1 0 904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_740
timestamp 1681620392
transform 1 0 912 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_208
timestamp 1681620392
transform 1 0 920 0 -1 1370
box -9 -3 26 105
use FILL  FILL_741
timestamp 1681620392
transform 1 0 936 0 -1 1370
box -8 -3 16 105
use FILL  FILL_742
timestamp 1681620392
transform 1 0 944 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_49
timestamp 1681620392
transform -1 0 992 0 -1 1370
box -8 -3 46 105
use FILL  FILL_743
timestamp 1681620392
transform 1 0 992 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_182
timestamp 1681620392
transform 1 0 1000 0 -1 1370
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_180
timestamp 1681620392
transform 1 0 1032 0 -1 1370
box -8 -3 104 105
use BUFX2  BUFX2_31
timestamp 1681620392
transform -1 0 1152 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_32
timestamp 1681620392
transform 1 0 1152 0 -1 1370
box -5 -3 28 105
use FILL  FILL_745
timestamp 1681620392
transform 1 0 1176 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_183
timestamp 1681620392
transform 1 0 1184 0 -1 1370
box -8 -3 34 105
use FILL  FILL_748
timestamp 1681620392
transform 1 0 1216 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_184
timestamp 1681620392
transform -1 0 1256 0 -1 1370
box -8 -3 34 105
use FILL  FILL_749
timestamp 1681620392
transform 1 0 1256 0 -1 1370
box -8 -3 16 105
use FILL  FILL_753
timestamp 1681620392
transform 1 0 1264 0 -1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_191
timestamp 1681620392
transform -1 0 1296 0 -1 1370
box -8 -3 32 105
use FILL  FILL_754
timestamp 1681620392
transform 1 0 1296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_755
timestamp 1681620392
transform 1 0 1304 0 -1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_72
timestamp 1681620392
transform 1 0 1312 0 -1 1370
box -8 -3 40 105
use FILL  FILL_756
timestamp 1681620392
transform 1 0 1344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_757
timestamp 1681620392
transform 1 0 1352 0 -1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_73
timestamp 1681620392
transform 1 0 1360 0 -1 1370
box -8 -3 40 105
use FILL  FILL_758
timestamp 1681620392
transform 1 0 1392 0 -1 1370
box -8 -3 16 105
use FILL  FILL_760
timestamp 1681620392
transform 1 0 1400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_782
timestamp 1681620392
transform 1 0 1408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_783
timestamp 1681620392
transform 1 0 1416 0 -1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_199
timestamp 1681620392
transform 1 0 1424 0 -1 1370
box -8 -3 32 105
use OAI21X1  OAI21X1_191
timestamp 1681620392
transform 1 0 1448 0 -1 1370
box -8 -3 34 105
use FILL  FILL_784
timestamp 1681620392
transform 1 0 1480 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_192
timestamp 1681620392
transform 1 0 1488 0 -1 1370
box -8 -3 34 105
use INVX2  INVX2_216
timestamp 1681620392
transform -1 0 1536 0 -1 1370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_187
timestamp 1681620392
transform 1 0 1536 0 -1 1370
box -8 -3 104 105
use INVX2  INVX2_217
timestamp 1681620392
transform 1 0 1632 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_218
timestamp 1681620392
transform 1 0 1648 0 -1 1370
box -9 -3 26 105
use OAI21X1  OAI21X1_193
timestamp 1681620392
transform 1 0 1664 0 -1 1370
box -8 -3 34 105
use NAND2X1  NAND2X1_200
timestamp 1681620392
transform -1 0 1720 0 -1 1370
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_188
timestamp 1681620392
transform 1 0 1720 0 -1 1370
box -8 -3 104 105
use INVX2  INVX2_219
timestamp 1681620392
transform 1 0 1816 0 -1 1370
box -9 -3 26 105
use OAI22X1  OAI22X1_52
timestamp 1681620392
transform -1 0 1872 0 -1 1370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_189
timestamp 1681620392
transform 1 0 1872 0 -1 1370
box -8 -3 104 105
use NAND2X1  NAND2X1_201
timestamp 1681620392
transform -1 0 1992 0 -1 1370
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_190
timestamp 1681620392
transform 1 0 1992 0 -1 1370
box -8 -3 104 105
use OAI22X1  OAI22X1_53
timestamp 1681620392
transform 1 0 2088 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_54
timestamp 1681620392
transform -1 0 2168 0 -1 1370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_191
timestamp 1681620392
transform 1 0 2168 0 -1 1370
box -8 -3 104 105
use NAND2X1  NAND2X1_202
timestamp 1681620392
transform 1 0 2264 0 -1 1370
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_192
timestamp 1681620392
transform 1 0 2288 0 -1 1370
box -8 -3 104 105
use INVX2  INVX2_220
timestamp 1681620392
transform 1 0 2384 0 -1 1370
box -9 -3 26 105
use OAI21X1  OAI21X1_194
timestamp 1681620392
transform 1 0 2400 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_195
timestamp 1681620392
transform -1 0 2464 0 -1 1370
box -8 -3 34 105
use INVX2  INVX2_221
timestamp 1681620392
transform 1 0 2464 0 -1 1370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_193
timestamp 1681620392
transform 1 0 2480 0 -1 1370
box -8 -3 104 105
use OAI22X1  OAI22X1_55
timestamp 1681620392
transform -1 0 2616 0 -1 1370
box -8 -3 46 105
use OAI21X1  OAI21X1_196
timestamp 1681620392
transform -1 0 2648 0 -1 1370
box -8 -3 34 105
use OAI22X1  OAI22X1_56
timestamp 1681620392
transform -1 0 2688 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_57
timestamp 1681620392
transform 1 0 2688 0 -1 1370
box -8 -3 46 105
use NAND2X1  NAND2X1_203
timestamp 1681620392
transform 1 0 2728 0 -1 1370
box -8 -3 32 105
use M3_M2  M3_M2_2862
timestamp 1681620392
transform 1 0 2780 0 1 1275
box -3 -3 3 3
use OAI21X1  OAI21X1_197
timestamp 1681620392
transform 1 0 2752 0 -1 1370
box -8 -3 34 105
use NAND2X1  NAND2X1_205
timestamp 1681620392
transform 1 0 2784 0 -1 1370
box -8 -3 32 105
use FILL  FILL_788
timestamp 1681620392
transform 1 0 2808 0 -1 1370
box -8 -3 16 105
use FILL  FILL_790
timestamp 1681620392
transform 1 0 2816 0 -1 1370
box -8 -3 16 105
use FILL  FILL_792
timestamp 1681620392
transform 1 0 2824 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_58
timestamp 1681620392
transform 1 0 2832 0 -1 1370
box -8 -3 46 105
use FILL  FILL_795
timestamp 1681620392
transform 1 0 2872 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_2863
timestamp 1681620392
transform 1 0 2892 0 1 1275
box -3 -3 3 3
use FILL  FILL_797
timestamp 1681620392
transform 1 0 2880 0 -1 1370
box -8 -3 16 105
use FILL  FILL_799
timestamp 1681620392
transform 1 0 2888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_801
timestamp 1681620392
transform 1 0 2896 0 -1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_70
timestamp 1681620392
transform 1 0 2904 0 -1 1370
box -8 -3 32 105
use INVX2  INVX2_224
timestamp 1681620392
transform 1 0 2928 0 -1 1370
box -9 -3 26 105
use FILL  FILL_803
timestamp 1681620392
transform 1 0 2944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_805
timestamp 1681620392
transform 1 0 2952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_808
timestamp 1681620392
transform 1 0 2960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_809
timestamp 1681620392
transform 1 0 2968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_810
timestamp 1681620392
transform 1 0 2976 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_225
timestamp 1681620392
transform 1 0 2984 0 -1 1370
box -9 -3 26 105
use FILL  FILL_811
timestamp 1681620392
transform 1 0 3000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_813
timestamp 1681620392
transform 1 0 3008 0 -1 1370
box -8 -3 16 105
use Project_Top_VIA0  Project_Top_VIA0_35
timestamp 1681620392
transform 1 0 3067 0 1 1270
box -10 -3 10 3
use M2_M1  M2_M1_3478
timestamp 1681620392
transform 1 0 84 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2889
timestamp 1681620392
transform 1 0 100 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_3349
timestamp 1681620392
transform 1 0 108 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_3360
timestamp 1681620392
transform 1 0 100 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_2899
timestamp 1681620392
transform 1 0 124 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_3361
timestamp 1681620392
transform 1 0 124 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_2926
timestamp 1681620392
transform 1 0 132 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2864
timestamp 1681620392
transform 1 0 164 0 1 1265
box -3 -3 3 3
use M2_M1  M2_M1_3362
timestamp 1681620392
transform 1 0 148 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3395
timestamp 1681620392
transform 1 0 132 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2872
timestamp 1681620392
transform 1 0 172 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2890
timestamp 1681620392
transform 1 0 180 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2927
timestamp 1681620392
transform 1 0 172 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_3396
timestamp 1681620392
transform 1 0 164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3479
timestamp 1681620392
transform 1 0 156 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3480
timestamp 1681620392
transform 1 0 172 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2873
timestamp 1681620392
transform 1 0 220 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2891
timestamp 1681620392
transform 1 0 220 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2900
timestamp 1681620392
transform 1 0 196 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2928
timestamp 1681620392
transform 1 0 188 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2959
timestamp 1681620392
transform 1 0 188 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_3350
timestamp 1681620392
transform 1 0 228 0 1 1235
box -2 -2 2 2
use M3_M2  M3_M2_2929
timestamp 1681620392
transform 1 0 212 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_3363
timestamp 1681620392
transform 1 0 220 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3397
timestamp 1681620392
transform 1 0 196 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3398
timestamp 1681620392
transform 1 0 212 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2874
timestamp 1681620392
transform 1 0 300 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_3351
timestamp 1681620392
transform 1 0 268 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_3364
timestamp 1681620392
transform 1 0 244 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3365
timestamp 1681620392
transform 1 0 252 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_2960
timestamp 1681620392
transform 1 0 244 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2901
timestamp 1681620392
transform 1 0 276 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_3366
timestamp 1681620392
transform 1 0 276 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_2930
timestamp 1681620392
transform 1 0 284 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2875
timestamp 1681620392
transform 1 0 332 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2892
timestamp 1681620392
transform 1 0 324 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2931
timestamp 1681620392
transform 1 0 316 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_3399
timestamp 1681620392
transform 1 0 260 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3400
timestamp 1681620392
transform 1 0 284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3401
timestamp 1681620392
transform 1 0 300 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2976
timestamp 1681620392
transform 1 0 244 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_3481
timestamp 1681620392
transform 1 0 308 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3482
timestamp 1681620392
transform 1 0 316 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2893
timestamp 1681620392
transform 1 0 348 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_3352
timestamp 1681620392
transform 1 0 356 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_3367
timestamp 1681620392
transform 1 0 332 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3368
timestamp 1681620392
transform 1 0 340 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3369
timestamp 1681620392
transform 1 0 348 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_2932
timestamp 1681620392
transform 1 0 356 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2902
timestamp 1681620392
transform 1 0 380 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_3370
timestamp 1681620392
transform 1 0 364 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3402
timestamp 1681620392
transform 1 0 332 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3403
timestamp 1681620392
transform 1 0 348 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2961
timestamp 1681620392
transform 1 0 356 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_3404
timestamp 1681620392
transform 1 0 372 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3483
timestamp 1681620392
transform 1 0 372 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2876
timestamp 1681620392
transform 1 0 412 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2894
timestamp 1681620392
transform 1 0 420 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_3353
timestamp 1681620392
transform 1 0 412 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_3354
timestamp 1681620392
transform 1 0 420 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_3371
timestamp 1681620392
transform 1 0 396 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3372
timestamp 1681620392
transform 1 0 404 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_2933
timestamp 1681620392
transform 1 0 420 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_3373
timestamp 1681620392
transform 1 0 428 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_2962
timestamp 1681620392
transform 1 0 396 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2963
timestamp 1681620392
transform 1 0 412 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_3484
timestamp 1681620392
transform 1 0 396 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2990
timestamp 1681620392
transform 1 0 396 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2877
timestamp 1681620392
transform 1 0 444 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2964
timestamp 1681620392
transform 1 0 436 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2903
timestamp 1681620392
transform 1 0 452 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2865
timestamp 1681620392
transform 1 0 492 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2878
timestamp 1681620392
transform 1 0 484 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_3355
timestamp 1681620392
transform 1 0 468 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_3374
timestamp 1681620392
transform 1 0 452 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_2977
timestamp 1681620392
transform 1 0 444 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2904
timestamp 1681620392
transform 1 0 476 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_3375
timestamp 1681620392
transform 1 0 492 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_2934
timestamp 1681620392
transform 1 0 500 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_3376
timestamp 1681620392
transform 1 0 508 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_2965
timestamp 1681620392
transform 1 0 492 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_3485
timestamp 1681620392
transform 1 0 484 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2966
timestamp 1681620392
transform 1 0 516 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2935
timestamp 1681620392
transform 1 0 532 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_3486
timestamp 1681620392
transform 1 0 524 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3487
timestamp 1681620392
transform 1 0 532 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3377
timestamp 1681620392
transform 1 0 572 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3405
timestamp 1681620392
transform 1 0 556 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2866
timestamp 1681620392
transform 1 0 612 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2867
timestamp 1681620392
transform 1 0 708 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2905
timestamp 1681620392
transform 1 0 700 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2936
timestamp 1681620392
transform 1 0 668 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_3406
timestamp 1681620392
transform 1 0 596 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3407
timestamp 1681620392
transform 1 0 612 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3408
timestamp 1681620392
transform 1 0 668 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3488
timestamp 1681620392
transform 1 0 580 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3489
timestamp 1681620392
transform 1 0 604 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3490
timestamp 1681620392
transform 1 0 692 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2991
timestamp 1681620392
transform 1 0 644 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2992
timestamp 1681620392
transform 1 0 692 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2937
timestamp 1681620392
transform 1 0 740 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_3409
timestamp 1681620392
transform 1 0 764 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3491
timestamp 1681620392
transform 1 0 716 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2993
timestamp 1681620392
transform 1 0 716 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2994
timestamp 1681620392
transform 1 0 764 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2895
timestamp 1681620392
transform 1 0 820 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2938
timestamp 1681620392
transform 1 0 820 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2906
timestamp 1681620392
transform 1 0 868 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_3378
timestamp 1681620392
transform 1 0 860 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3410
timestamp 1681620392
transform 1 0 812 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3411
timestamp 1681620392
transform 1 0 844 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2896
timestamp 1681620392
transform 1 0 988 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2907
timestamp 1681620392
transform 1 0 980 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2939
timestamp 1681620392
transform 1 0 884 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2940
timestamp 1681620392
transform 1 0 972 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_3412
timestamp 1681620392
transform 1 0 876 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3413
timestamp 1681620392
transform 1 0 884 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3414
timestamp 1681620392
transform 1 0 924 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3492
timestamp 1681620392
transform 1 0 820 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3493
timestamp 1681620392
transform 1 0 836 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3494
timestamp 1681620392
transform 1 0 852 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3495
timestamp 1681620392
transform 1 0 860 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2995
timestamp 1681620392
transform 1 0 836 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2996
timestamp 1681620392
transform 1 0 860 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_3496
timestamp 1681620392
transform 1 0 900 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2997
timestamp 1681620392
transform 1 0 924 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3021
timestamp 1681620392
transform 1 0 900 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2941
timestamp 1681620392
transform 1 0 1036 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2942
timestamp 1681620392
transform 1 0 1084 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_3415
timestamp 1681620392
transform 1 0 996 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3416
timestamp 1681620392
transform 1 0 1036 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3497
timestamp 1681620392
transform 1 0 1012 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_3022
timestamp 1681620392
transform 1 0 1012 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3023
timestamp 1681620392
transform 1 0 1076 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2908
timestamp 1681620392
transform 1 0 1108 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_3417
timestamp 1681620392
transform 1 0 1108 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3418
timestamp 1681620392
transform 1 0 1116 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2943
timestamp 1681620392
transform 1 0 1132 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_3419
timestamp 1681620392
transform 1 0 1132 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3498
timestamp 1681620392
transform 1 0 1124 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3548
timestamp 1681620392
transform 1 0 1132 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_3024
timestamp 1681620392
transform 1 0 1132 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2909
timestamp 1681620392
transform 1 0 1164 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2944
timestamp 1681620392
transform 1 0 1156 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2945
timestamp 1681620392
transform 1 0 1196 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_3420
timestamp 1681620392
transform 1 0 1156 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3421
timestamp 1681620392
transform 1 0 1220 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3499
timestamp 1681620392
transform 1 0 1156 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3500
timestamp 1681620392
transform 1 0 1172 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2998
timestamp 1681620392
transform 1 0 1220 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3025
timestamp 1681620392
transform 1 0 1252 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2910
timestamp 1681620392
transform 1 0 1292 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2946
timestamp 1681620392
transform 1 0 1268 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2947
timestamp 1681620392
transform 1 0 1284 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_3422
timestamp 1681620392
transform 1 0 1268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3423
timestamp 1681620392
transform 1 0 1276 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2978
timestamp 1681620392
transform 1 0 1276 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_3424
timestamp 1681620392
transform 1 0 1284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3425
timestamp 1681620392
transform 1 0 1300 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3426
timestamp 1681620392
transform 1 0 1316 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3501
timestamp 1681620392
transform 1 0 1284 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3502
timestamp 1681620392
transform 1 0 1292 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3503
timestamp 1681620392
transform 1 0 1308 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2999
timestamp 1681620392
transform 1 0 1308 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3026
timestamp 1681620392
transform 1 0 1284 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_3379
timestamp 1681620392
transform 1 0 1332 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3504
timestamp 1681620392
transform 1 0 1332 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3356
timestamp 1681620392
transform 1 0 1364 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_3380
timestamp 1681620392
transform 1 0 1364 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3427
timestamp 1681620392
transform 1 0 1356 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3428
timestamp 1681620392
transform 1 0 1372 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2979
timestamp 1681620392
transform 1 0 1364 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_3381
timestamp 1681620392
transform 1 0 1388 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_2911
timestamp 1681620392
transform 1 0 1500 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2912
timestamp 1681620392
transform 1 0 1604 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_3429
timestamp 1681620392
transform 1 0 1404 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3430
timestamp 1681620392
transform 1 0 1412 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3431
timestamp 1681620392
transform 1 0 1452 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3432
timestamp 1681620392
transform 1 0 1508 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3433
timestamp 1681620392
transform 1 0 1572 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3434
timestamp 1681620392
transform 1 0 1604 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3505
timestamp 1681620392
transform 1 0 1380 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3506
timestamp 1681620392
transform 1 0 1388 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2980
timestamp 1681620392
transform 1 0 1396 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_3000
timestamp 1681620392
transform 1 0 1388 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_3507
timestamp 1681620392
transform 1 0 1428 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_3001
timestamp 1681620392
transform 1 0 1452 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_3508
timestamp 1681620392
transform 1 0 1524 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2981
timestamp 1681620392
transform 1 0 1572 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2982
timestamp 1681620392
transform 1 0 1596 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_3549
timestamp 1681620392
transform 1 0 1612 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_3027
timestamp 1681620392
transform 1 0 1524 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_3357
timestamp 1681620392
transform 1 0 1644 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_3358
timestamp 1681620392
transform 1 0 1652 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_3382
timestamp 1681620392
transform 1 0 1636 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3383
timestamp 1681620392
transform 1 0 1660 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3435
timestamp 1681620392
transform 1 0 1628 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3436
timestamp 1681620392
transform 1 0 1652 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3509
timestamp 1681620392
transform 1 0 1628 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2983
timestamp 1681620392
transform 1 0 1652 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_3002
timestamp 1681620392
transform 1 0 1628 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3003
timestamp 1681620392
transform 1 0 1644 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2913
timestamp 1681620392
transform 1 0 1676 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_3384
timestamp 1681620392
transform 1 0 1676 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3359
timestamp 1681620392
transform 1 0 1700 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_3385
timestamp 1681620392
transform 1 0 1708 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3437
timestamp 1681620392
transform 1 0 1692 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2914
timestamp 1681620392
transform 1 0 1852 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2948
timestamp 1681620392
transform 1 0 1828 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2949
timestamp 1681620392
transform 1 0 1900 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_3438
timestamp 1681620392
transform 1 0 1724 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3439
timestamp 1681620392
transform 1 0 1732 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3440
timestamp 1681620392
transform 1 0 1764 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3441
timestamp 1681620392
transform 1 0 1828 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3510
timestamp 1681620392
transform 1 0 1716 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_3004
timestamp 1681620392
transform 1 0 1692 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2984
timestamp 1681620392
transform 1 0 1724 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2967
timestamp 1681620392
transform 1 0 1836 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_3442
timestamp 1681620392
transform 1 0 1852 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2968
timestamp 1681620392
transform 1 0 1868 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_3443
timestamp 1681620392
transform 1 0 1876 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3444
timestamp 1681620392
transform 1 0 1892 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3445
timestamp 1681620392
transform 1 0 1900 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2969
timestamp 1681620392
transform 1 0 1908 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2868
timestamp 1681620392
transform 1 0 1988 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2897
timestamp 1681620392
transform 1 0 2036 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_3386
timestamp 1681620392
transform 1 0 1932 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_2950
timestamp 1681620392
transform 1 0 1972 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2951
timestamp 1681620392
transform 1 0 1988 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2915
timestamp 1681620392
transform 1 0 2116 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2952
timestamp 1681620392
transform 1 0 2092 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_3446
timestamp 1681620392
transform 1 0 1932 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3447
timestamp 1681620392
transform 1 0 1972 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3448
timestamp 1681620392
transform 1 0 2028 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3449
timestamp 1681620392
transform 1 0 2092 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3511
timestamp 1681620392
transform 1 0 1812 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3512
timestamp 1681620392
transform 1 0 1828 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3513
timestamp 1681620392
transform 1 0 1844 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3514
timestamp 1681620392
transform 1 0 1860 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3515
timestamp 1681620392
transform 1 0 1868 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3516
timestamp 1681620392
transform 1 0 1884 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3517
timestamp 1681620392
transform 1 0 1900 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3518
timestamp 1681620392
transform 1 0 1908 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_3005
timestamp 1681620392
transform 1 0 1828 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3028
timestamp 1681620392
transform 1 0 1812 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3006
timestamp 1681620392
transform 1 0 1892 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2985
timestamp 1681620392
transform 1 0 1924 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_3519
timestamp 1681620392
transform 1 0 1948 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_3007
timestamp 1681620392
transform 1 0 1916 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3008
timestamp 1681620392
transform 1 0 1932 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3029
timestamp 1681620392
transform 1 0 1908 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_3520
timestamp 1681620392
transform 1 0 2044 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2986
timestamp 1681620392
transform 1 0 2068 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_3030
timestamp 1681620392
transform 1 0 2028 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2953
timestamp 1681620392
transform 1 0 2148 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2898
timestamp 1681620392
transform 1 0 2228 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2916
timestamp 1681620392
transform 1 0 2172 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_3387
timestamp 1681620392
transform 1 0 2172 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3450
timestamp 1681620392
transform 1 0 2156 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3521
timestamp 1681620392
transform 1 0 2148 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2987
timestamp 1681620392
transform 1 0 2156 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2917
timestamp 1681620392
transform 1 0 2284 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_3388
timestamp 1681620392
transform 1 0 2276 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3451
timestamp 1681620392
transform 1 0 2212 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3452
timestamp 1681620392
transform 1 0 2276 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3453
timestamp 1681620392
transform 1 0 2284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3522
timestamp 1681620392
transform 1 0 2172 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3523
timestamp 1681620392
transform 1 0 2188 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_3009
timestamp 1681620392
transform 1 0 2132 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3010
timestamp 1681620392
transform 1 0 2148 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3011
timestamp 1681620392
transform 1 0 2172 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3012
timestamp 1681620392
transform 1 0 2212 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2869
timestamp 1681620392
transform 1 0 2356 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2879
timestamp 1681620392
transform 1 0 2348 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2918
timestamp 1681620392
transform 1 0 2316 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2919
timestamp 1681620392
transform 1 0 2332 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_3389
timestamp 1681620392
transform 1 0 2316 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3454
timestamp 1681620392
transform 1 0 2308 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3455
timestamp 1681620392
transform 1 0 2316 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3524
timestamp 1681620392
transform 1 0 2292 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3525
timestamp 1681620392
transform 1 0 2300 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_3031
timestamp 1681620392
transform 1 0 2300 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2920
timestamp 1681620392
transform 1 0 2364 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2870
timestamp 1681620392
transform 1 0 2396 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2880
timestamp 1681620392
transform 1 0 2396 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2881
timestamp 1681620392
transform 1 0 2444 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2882
timestamp 1681620392
transform 1 0 2460 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_3390
timestamp 1681620392
transform 1 0 2372 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3456
timestamp 1681620392
transform 1 0 2340 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3457
timestamp 1681620392
transform 1 0 2348 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3458
timestamp 1681620392
transform 1 0 2356 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3459
timestamp 1681620392
transform 1 0 2364 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3526
timestamp 1681620392
transform 1 0 2324 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2883
timestamp 1681620392
transform 1 0 2492 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2921
timestamp 1681620392
transform 1 0 2476 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_3391
timestamp 1681620392
transform 1 0 2476 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3460
timestamp 1681620392
transform 1 0 2436 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3461
timestamp 1681620392
transform 1 0 2468 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2884
timestamp 1681620392
transform 1 0 2524 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2885
timestamp 1681620392
transform 1 0 2572 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2922
timestamp 1681620392
transform 1 0 2588 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2954
timestamp 1681620392
transform 1 0 2500 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2955
timestamp 1681620392
transform 1 0 2596 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_3462
timestamp 1681620392
transform 1 0 2492 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3463
timestamp 1681620392
transform 1 0 2500 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3464
timestamp 1681620392
transform 1 0 2540 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3465
timestamp 1681620392
transform 1 0 2596 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3466
timestamp 1681620392
transform 1 0 2604 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3527
timestamp 1681620392
transform 1 0 2388 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3528
timestamp 1681620392
transform 1 0 2476 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_3013
timestamp 1681620392
transform 1 0 2388 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3014
timestamp 1681620392
transform 1 0 2420 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3015
timestamp 1681620392
transform 1 0 2476 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3032
timestamp 1681620392
transform 1 0 2452 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_3529
timestamp 1681620392
transform 1 0 2516 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_3016
timestamp 1681620392
transform 1 0 2540 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3017
timestamp 1681620392
transform 1 0 2596 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3033
timestamp 1681620392
transform 1 0 2532 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2886
timestamp 1681620392
transform 1 0 2620 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2923
timestamp 1681620392
transform 1 0 2612 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_3467
timestamp 1681620392
transform 1 0 2612 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3530
timestamp 1681620392
transform 1 0 2612 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2956
timestamp 1681620392
transform 1 0 2628 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_3468
timestamp 1681620392
transform 1 0 2636 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3531
timestamp 1681620392
transform 1 0 2628 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2970
timestamp 1681620392
transform 1 0 2644 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_3532
timestamp 1681620392
transform 1 0 2644 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3392
timestamp 1681620392
transform 1 0 2668 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_2871
timestamp 1681620392
transform 1 0 2684 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2971
timestamp 1681620392
transform 1 0 2676 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_3469
timestamp 1681620392
transform 1 0 2684 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2988
timestamp 1681620392
transform 1 0 2684 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_3533
timestamp 1681620392
transform 1 0 2692 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_2887
timestamp 1681620392
transform 1 0 2708 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2972
timestamp 1681620392
transform 1 0 2716 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_3534
timestamp 1681620392
transform 1 0 2708 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_3034
timestamp 1681620392
transform 1 0 2700 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2888
timestamp 1681620392
transform 1 0 2740 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2924
timestamp 1681620392
transform 1 0 2772 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2925
timestamp 1681620392
transform 1 0 2788 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2957
timestamp 1681620392
transform 1 0 2740 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2958
timestamp 1681620392
transform 1 0 2764 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_3393
timestamp 1681620392
transform 1 0 2788 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3470
timestamp 1681620392
transform 1 0 2748 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2973
timestamp 1681620392
transform 1 0 2756 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_3471
timestamp 1681620392
transform 1 0 2764 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3535
timestamp 1681620392
transform 1 0 2740 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3536
timestamp 1681620392
transform 1 0 2756 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3537
timestamp 1681620392
transform 1 0 2764 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_3018
timestamp 1681620392
transform 1 0 2756 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2974
timestamp 1681620392
transform 1 0 2788 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_3472
timestamp 1681620392
transform 1 0 2812 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_2975
timestamp 1681620392
transform 1 0 2820 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_3473
timestamp 1681620392
transform 1 0 2836 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3538
timestamp 1681620392
transform 1 0 2796 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3539
timestamp 1681620392
transform 1 0 2804 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3540
timestamp 1681620392
transform 1 0 2812 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3541
timestamp 1681620392
transform 1 0 2820 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3550
timestamp 1681620392
transform 1 0 2796 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_2989
timestamp 1681620392
transform 1 0 2836 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_3542
timestamp 1681620392
transform 1 0 2844 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_3035
timestamp 1681620392
transform 1 0 2796 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3036
timestamp 1681620392
transform 1 0 2820 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_3543
timestamp 1681620392
transform 1 0 2868 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3394
timestamp 1681620392
transform 1 0 2908 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3474
timestamp 1681620392
transform 1 0 2884 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3475
timestamp 1681620392
transform 1 0 2892 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3476
timestamp 1681620392
transform 1 0 2924 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3477
timestamp 1681620392
transform 1 0 2940 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3544
timestamp 1681620392
transform 1 0 2908 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3545
timestamp 1681620392
transform 1 0 2916 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3546
timestamp 1681620392
transform 1 0 2932 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3547
timestamp 1681620392
transform 1 0 2948 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_3019
timestamp 1681620392
transform 1 0 2908 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3020
timestamp 1681620392
transform 1 0 2948 0 1 1195
box -3 -3 3 3
use Project_Top_VIA0  Project_Top_VIA0_36
timestamp 1681620392
transform 1 0 48 0 1 1170
box -10 -3 10 3
use FILL  FILL_814
timestamp 1681620392
transform 1 0 72 0 1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_207
timestamp 1681620392
transform 1 0 80 0 1 1170
box -8 -3 32 105
use FILL  FILL_815
timestamp 1681620392
transform 1 0 104 0 1 1170
box -8 -3 16 105
use FILL  FILL_816
timestamp 1681620392
transform 1 0 112 0 1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_74
timestamp 1681620392
transform 1 0 120 0 1 1170
box -8 -3 40 105
use INVX2  INVX2_226
timestamp 1681620392
transform 1 0 152 0 1 1170
box -9 -3 26 105
use FILL  FILL_817
timestamp 1681620392
transform 1 0 168 0 1 1170
box -8 -3 16 105
use FILL  FILL_819
timestamp 1681620392
transform 1 0 176 0 1 1170
box -8 -3 16 105
use AND2X2  AND2X2_20
timestamp 1681620392
transform 1 0 184 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_75
timestamp 1681620392
transform -1 0 248 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_76
timestamp 1681620392
transform 1 0 248 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_21
timestamp 1681620392
transform -1 0 312 0 1 1170
box -8 -3 40 105
use NAND2X1  NAND2X1_208
timestamp 1681620392
transform 1 0 312 0 1 1170
box -8 -3 32 105
use NAND3X1  NAND3X1_77
timestamp 1681620392
transform 1 0 336 0 1 1170
box -8 -3 40 105
use OAI21X1  OAI21X1_200
timestamp 1681620392
transform 1 0 368 0 1 1170
box -8 -3 34 105
use NAND3X1  NAND3X1_78
timestamp 1681620392
transform -1 0 432 0 1 1170
box -8 -3 40 105
use FILL  FILL_821
timestamp 1681620392
transform 1 0 432 0 1 1170
box -8 -3 16 105
use FILL  FILL_822
timestamp 1681620392
transform 1 0 440 0 1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_79
timestamp 1681620392
transform 1 0 448 0 1 1170
box -8 -3 40 105
use FILL  FILL_823
timestamp 1681620392
transform 1 0 480 0 1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_209
timestamp 1681620392
transform 1 0 488 0 1 1170
box -8 -3 32 105
use FILL  FILL_824
timestamp 1681620392
transform 1 0 512 0 1 1170
box -8 -3 16 105
use FILL  FILL_825
timestamp 1681620392
transform 1 0 520 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_227
timestamp 1681620392
transform 1 0 528 0 1 1170
box -9 -3 26 105
use OAI21X1  OAI21X1_201
timestamp 1681620392
transform 1 0 544 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_202
timestamp 1681620392
transform -1 0 608 0 1 1170
box -8 -3 34 105
use M3_M2  M3_M2_3037
timestamp 1681620392
transform 1 0 636 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3038
timestamp 1681620392
transform 1 0 652 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_195
timestamp 1681620392
transform -1 0 704 0 1 1170
box -8 -3 104 105
use M3_M2  M3_M2_3039
timestamp 1681620392
transform 1 0 724 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3040
timestamp 1681620392
transform 1 0 756 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_196
timestamp 1681620392
transform 1 0 704 0 1 1170
box -8 -3 104 105
use M3_M2  M3_M2_3041
timestamp 1681620392
transform 1 0 820 0 1 1175
box -3 -3 3 3
use INVX2  INVX2_228
timestamp 1681620392
transform 1 0 800 0 1 1170
box -9 -3 26 105
use OAI22X1  OAI22X1_59
timestamp 1681620392
transform 1 0 816 0 1 1170
box -8 -3 46 105
use M3_M2  M3_M2_3042
timestamp 1681620392
transform 1 0 876 0 1 1175
box -3 -3 3 3
use OAI21X1  OAI21X1_203
timestamp 1681620392
transform -1 0 888 0 1 1170
box -8 -3 34 105
use M3_M2  M3_M2_3043
timestamp 1681620392
transform 1 0 908 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_197
timestamp 1681620392
transform 1 0 888 0 1 1170
box -8 -3 104 105
use M3_M2  M3_M2_3044
timestamp 1681620392
transform 1 0 996 0 1 1175
box -3 -3 3 3
use INVX2  INVX2_229
timestamp 1681620392
transform 1 0 984 0 1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_198
timestamp 1681620392
transform 1 0 1000 0 1 1170
box -8 -3 104 105
use INVX2  INVX2_230
timestamp 1681620392
transform 1 0 1096 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_231
timestamp 1681620392
transform -1 0 1128 0 1 1170
box -9 -3 26 105
use AOI21X1  AOI21X1_21
timestamp 1681620392
transform -1 0 1160 0 1 1170
box -7 -3 39 105
use M3_M2  M3_M2_3045
timestamp 1681620392
transform 1 0 1204 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_199
timestamp 1681620392
transform 1 0 1160 0 1 1170
box -8 -3 104 105
use INVX2  INVX2_232
timestamp 1681620392
transform 1 0 1256 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_233
timestamp 1681620392
transform -1 0 1288 0 1 1170
box -9 -3 26 105
use OAI22X1  OAI22X1_60
timestamp 1681620392
transform 1 0 1288 0 1 1170
box -8 -3 46 105
use FILL  FILL_826
timestamp 1681620392
transform 1 0 1328 0 1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_80
timestamp 1681620392
transform -1 0 1368 0 1 1170
box -8 -3 40 105
use INVX2  INVX2_234
timestamp 1681620392
transform -1 0 1384 0 1 1170
box -9 -3 26 105
use OAI21X1  OAI21X1_204
timestamp 1681620392
transform -1 0 1416 0 1 1170
box -8 -3 34 105
use M3_M2  M3_M2_3046
timestamp 1681620392
transform 1 0 1444 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_200
timestamp 1681620392
transform 1 0 1416 0 1 1170
box -8 -3 104 105
use M3_M2  M3_M2_3047
timestamp 1681620392
transform 1 0 1532 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3048
timestamp 1681620392
transform 1 0 1588 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_201
timestamp 1681620392
transform 1 0 1512 0 1 1170
box -8 -3 104 105
use NOR2X1  NOR2X1_71
timestamp 1681620392
transform 1 0 1608 0 1 1170
box -8 -3 32 105
use NAND3X1  NAND3X1_81
timestamp 1681620392
transform -1 0 1664 0 1 1170
box -8 -3 40 105
use FILL  FILL_827
timestamp 1681620392
transform 1 0 1664 0 1 1170
box -8 -3 16 105
use FILL  FILL_828
timestamp 1681620392
transform 1 0 1672 0 1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_82
timestamp 1681620392
transform 1 0 1680 0 1 1170
box -8 -3 40 105
use INVX2  INVX2_235
timestamp 1681620392
transform 1 0 1712 0 1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_202
timestamp 1681620392
transform -1 0 1824 0 1 1170
box -8 -3 104 105
use OAI22X1  OAI22X1_61
timestamp 1681620392
transform 1 0 1824 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_62
timestamp 1681620392
transform -1 0 1904 0 1 1170
box -8 -3 46 105
use OAI21X1  OAI21X1_205
timestamp 1681620392
transform 1 0 1904 0 1 1170
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_203
timestamp 1681620392
transform 1 0 1936 0 1 1170
box -8 -3 104 105
use M3_M2  M3_M2_3049
timestamp 1681620392
transform 1 0 2108 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_204
timestamp 1681620392
transform 1 0 2032 0 1 1170
box -8 -3 104 105
use M3_M2  M3_M2_3050
timestamp 1681620392
transform 1 0 2140 0 1 1175
box -3 -3 3 3
use INVX2  INVX2_236
timestamp 1681620392
transform 1 0 2128 0 1 1170
box -9 -3 26 105
use OAI21X1  OAI21X1_206
timestamp 1681620392
transform 1 0 2144 0 1 1170
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_205
timestamp 1681620392
transform 1 0 2176 0 1 1170
box -8 -3 104 105
use NAND2X1  NAND2X1_210
timestamp 1681620392
transform -1 0 2296 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_211
timestamp 1681620392
transform 1 0 2296 0 1 1170
box -8 -3 32 105
use OAI21X1  OAI21X1_207
timestamp 1681620392
transform -1 0 2352 0 1 1170
box -8 -3 34 105
use NAND2X1  NAND2X1_212
timestamp 1681620392
transform 1 0 2352 0 1 1170
box -8 -3 32 105
use M3_M2  M3_M2_3051
timestamp 1681620392
transform 1 0 2420 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_206
timestamp 1681620392
transform 1 0 2376 0 1 1170
box -8 -3 104 105
use OAI21X1  OAI21X1_208
timestamp 1681620392
transform -1 0 2504 0 1 1170
box -8 -3 34 105
use M3_M2  M3_M2_3052
timestamp 1681620392
transform 1 0 2516 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3053
timestamp 1681620392
transform 1 0 2556 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_207
timestamp 1681620392
transform 1 0 2504 0 1 1170
box -8 -3 104 105
use M3_M2  M3_M2_3054
timestamp 1681620392
transform 1 0 2620 0 1 1175
box -3 -3 3 3
use INVX2  INVX2_237
timestamp 1681620392
transform -1 0 2616 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_238
timestamp 1681620392
transform -1 0 2632 0 1 1170
box -9 -3 26 105
use FILL  FILL_829
timestamp 1681620392
transform 1 0 2632 0 1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_209
timestamp 1681620392
transform 1 0 2640 0 1 1170
box -8 -3 34 105
use FILL  FILL_830
timestamp 1681620392
transform 1 0 2672 0 1 1170
box -8 -3 16 105
use FILL  FILL_831
timestamp 1681620392
transform 1 0 2680 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_3055
timestamp 1681620392
transform 1 0 2700 0 1 1175
box -3 -3 3 3
use FILL  FILL_832
timestamp 1681620392
transform 1 0 2688 0 1 1170
box -8 -3 16 105
use FILL  FILL_833
timestamp 1681620392
transform 1 0 2696 0 1 1170
box -8 -3 16 105
use FILL  FILL_834
timestamp 1681620392
transform 1 0 2704 0 1 1170
box -8 -3 16 105
use FILL  FILL_893
timestamp 1681620392
transform 1 0 2712 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_68
timestamp 1681620392
transform 1 0 2720 0 1 1170
box -8 -3 46 105
use OAI21X1  OAI21X1_218
timestamp 1681620392
transform 1 0 2760 0 1 1170
box -8 -3 34 105
use NOR2X1  NOR2X1_74
timestamp 1681620392
transform 1 0 2792 0 1 1170
box -8 -3 32 105
use AOI22X1  AOI22X1_29
timestamp 1681620392
transform -1 0 2856 0 1 1170
box -8 -3 46 105
use FILL  FILL_894
timestamp 1681620392
transform 1 0 2856 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_3056
timestamp 1681620392
transform 1 0 2876 0 1 1175
box -3 -3 3 3
use FILL  FILL_895
timestamp 1681620392
transform 1 0 2864 0 1 1170
box -8 -3 16 105
use FILL  FILL_896
timestamp 1681620392
transform 1 0 2872 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_3057
timestamp 1681620392
transform 1 0 2916 0 1 1175
box -3 -3 3 3
use OAI21X1  OAI21X1_219
timestamp 1681620392
transform 1 0 2880 0 1 1170
box -8 -3 34 105
use OAI22X1  OAI22X1_69
timestamp 1681620392
transform 1 0 2912 0 1 1170
box -8 -3 46 105
use FILL  FILL_897
timestamp 1681620392
transform 1 0 2952 0 1 1170
box -8 -3 16 105
use FILL  FILL_911
timestamp 1681620392
transform 1 0 2960 0 1 1170
box -8 -3 16 105
use FILL  FILL_912
timestamp 1681620392
transform 1 0 2968 0 1 1170
box -8 -3 16 105
use FILL  FILL_913
timestamp 1681620392
transform 1 0 2976 0 1 1170
box -8 -3 16 105
use FILL  FILL_914
timestamp 1681620392
transform 1 0 2984 0 1 1170
box -8 -3 16 105
use FILL  FILL_915
timestamp 1681620392
transform 1 0 2992 0 1 1170
box -8 -3 16 105
use FILL  FILL_916
timestamp 1681620392
transform 1 0 3000 0 1 1170
box -8 -3 16 105
use FILL  FILL_919
timestamp 1681620392
transform 1 0 3008 0 1 1170
box -8 -3 16 105
use Project_Top_VIA0  Project_Top_VIA0_37
timestamp 1681620392
transform 1 0 3043 0 1 1170
box -10 -3 10 3
use M3_M2  M3_M2_3074
timestamp 1681620392
transform 1 0 164 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_3556
timestamp 1681620392
transform 1 0 84 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3633
timestamp 1681620392
transform 1 0 132 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3075
timestamp 1681620392
transform 1 0 180 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3089
timestamp 1681620392
transform 1 0 180 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3634
timestamp 1681620392
transform 1 0 180 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3714
timestamp 1681620392
transform 1 0 172 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_3058
timestamp 1681620392
transform 1 0 196 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3090
timestamp 1681620392
transform 1 0 220 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3557
timestamp 1681620392
transform 1 0 220 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3635
timestamp 1681620392
transform 1 0 196 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3136
timestamp 1681620392
transform 1 0 212 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_3715
timestamp 1681620392
transform 1 0 212 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3730
timestamp 1681620392
transform 1 0 204 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_3636
timestamp 1681620392
transform 1 0 236 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3059
timestamp 1681620392
transform 1 0 260 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_3551
timestamp 1681620392
transform 1 0 252 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_3091
timestamp 1681620392
transform 1 0 284 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3552
timestamp 1681620392
transform 1 0 292 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_3558
timestamp 1681620392
transform 1 0 300 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3559
timestamp 1681620392
transform 1 0 308 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3560
timestamp 1681620392
transform 1 0 324 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3637
timestamp 1681620392
transform 1 0 292 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3638
timestamp 1681620392
transform 1 0 316 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3155
timestamp 1681620392
transform 1 0 308 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3183
timestamp 1681620392
transform 1 0 300 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_3561
timestamp 1681620392
transform 1 0 340 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_3137
timestamp 1681620392
transform 1 0 340 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3184
timestamp 1681620392
transform 1 0 348 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3124
timestamp 1681620392
transform 1 0 372 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_3639
timestamp 1681620392
transform 1 0 372 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3076
timestamp 1681620392
transform 1 0 412 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3092
timestamp 1681620392
transform 1 0 396 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3093
timestamp 1681620392
transform 1 0 452 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3562
timestamp 1681620392
transform 1 0 396 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3563
timestamp 1681620392
transform 1 0 412 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_3125
timestamp 1681620392
transform 1 0 468 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_3077
timestamp 1681620392
transform 1 0 548 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3094
timestamp 1681620392
transform 1 0 548 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3564
timestamp 1681620392
transform 1 0 500 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3565
timestamp 1681620392
transform 1 0 516 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3566
timestamp 1681620392
transform 1 0 532 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3640
timestamp 1681620392
transform 1 0 388 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3641
timestamp 1681620392
transform 1 0 412 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3642
timestamp 1681620392
transform 1 0 420 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3643
timestamp 1681620392
transform 1 0 452 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3156
timestamp 1681620392
transform 1 0 388 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3157
timestamp 1681620392
transform 1 0 412 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3185
timestamp 1681620392
transform 1 0 500 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3215
timestamp 1681620392
transform 1 0 420 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3126
timestamp 1681620392
transform 1 0 540 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_3567
timestamp 1681620392
transform 1 0 548 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3644
timestamp 1681620392
transform 1 0 524 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3645
timestamp 1681620392
transform 1 0 540 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3646
timestamp 1681620392
transform 1 0 548 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3158
timestamp 1681620392
transform 1 0 524 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3159
timestamp 1681620392
transform 1 0 548 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_3716
timestamp 1681620392
transform 1 0 556 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_3186
timestamp 1681620392
transform 1 0 540 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3216
timestamp 1681620392
transform 1 0 516 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3078
timestamp 1681620392
transform 1 0 580 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3095
timestamp 1681620392
transform 1 0 580 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3568
timestamp 1681620392
transform 1 0 580 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_3138
timestamp 1681620392
transform 1 0 604 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_3569
timestamp 1681620392
transform 1 0 620 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3647
timestamp 1681620392
transform 1 0 612 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3187
timestamp 1681620392
transform 1 0 612 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3127
timestamp 1681620392
transform 1 0 628 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_3648
timestamp 1681620392
transform 1 0 628 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3204
timestamp 1681620392
transform 1 0 628 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_3717
timestamp 1681620392
transform 1 0 644 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_3096
timestamp 1681620392
transform 1 0 676 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3570
timestamp 1681620392
transform 1 0 652 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_3128
timestamp 1681620392
transform 1 0 660 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_3571
timestamp 1681620392
transform 1 0 676 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3649
timestamp 1681620392
transform 1 0 668 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3650
timestamp 1681620392
transform 1 0 676 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3160
timestamp 1681620392
transform 1 0 660 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3188
timestamp 1681620392
transform 1 0 676 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3060
timestamp 1681620392
transform 1 0 724 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3097
timestamp 1681620392
transform 1 0 748 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3572
timestamp 1681620392
transform 1 0 708 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3573
timestamp 1681620392
transform 1 0 724 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_3129
timestamp 1681620392
transform 1 0 748 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_3139
timestamp 1681620392
transform 1 0 724 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_3651
timestamp 1681620392
transform 1 0 748 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3652
timestamp 1681620392
transform 1 0 804 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3098
timestamp 1681620392
transform 1 0 820 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3574
timestamp 1681620392
transform 1 0 820 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3653
timestamp 1681620392
transform 1 0 828 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3161
timestamp 1681620392
transform 1 0 828 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_3575
timestamp 1681620392
transform 1 0 868 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3576
timestamp 1681620392
transform 1 0 876 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3654
timestamp 1681620392
transform 1 0 852 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3655
timestamp 1681620392
transform 1 0 868 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3577
timestamp 1681620392
transform 1 0 908 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3656
timestamp 1681620392
transform 1 0 900 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3657
timestamp 1681620392
transform 1 0 916 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3189
timestamp 1681620392
transform 1 0 876 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3162
timestamp 1681620392
transform 1 0 916 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3205
timestamp 1681620392
transform 1 0 908 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3163
timestamp 1681620392
transform 1 0 932 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3061
timestamp 1681620392
transform 1 0 948 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3062
timestamp 1681620392
transform 1 0 972 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3099
timestamp 1681620392
transform 1 0 1012 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3100
timestamp 1681620392
transform 1 0 1028 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3578
timestamp 1681620392
transform 1 0 948 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3658
timestamp 1681620392
transform 1 0 996 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3164
timestamp 1681620392
transform 1 0 996 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3079
timestamp 1681620392
transform 1 0 1052 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_3553
timestamp 1681620392
transform 1 0 1052 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_3579
timestamp 1681620392
transform 1 0 1068 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3659
timestamp 1681620392
transform 1 0 1044 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3660
timestamp 1681620392
transform 1 0 1052 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3140
timestamp 1681620392
transform 1 0 1068 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3063
timestamp 1681620392
transform 1 0 1092 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3064
timestamp 1681620392
transform 1 0 1172 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3101
timestamp 1681620392
transform 1 0 1092 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3580
timestamp 1681620392
transform 1 0 1092 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3661
timestamp 1681620392
transform 1 0 1076 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3165
timestamp 1681620392
transform 1 0 1052 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3141
timestamp 1681620392
transform 1 0 1116 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_3662
timestamp 1681620392
transform 1 0 1140 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3663
timestamp 1681620392
transform 1 0 1172 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3206
timestamp 1681620392
transform 1 0 1076 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3065
timestamp 1681620392
transform 1 0 1292 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3066
timestamp 1681620392
transform 1 0 1324 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_3554
timestamp 1681620392
transform 1 0 1220 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_3581
timestamp 1681620392
transform 1 0 1204 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3664
timestamp 1681620392
transform 1 0 1196 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3582
timestamp 1681620392
transform 1 0 1236 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3583
timestamp 1681620392
transform 1 0 1324 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3584
timestamp 1681620392
transform 1 0 1340 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3585
timestamp 1681620392
transform 1 0 1356 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3586
timestamp 1681620392
transform 1 0 1364 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3665
timestamp 1681620392
transform 1 0 1220 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3666
timestamp 1681620392
transform 1 0 1260 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3667
timestamp 1681620392
transform 1 0 1316 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3668
timestamp 1681620392
transform 1 0 1332 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3669
timestamp 1681620392
transform 1 0 1348 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3670
timestamp 1681620392
transform 1 0 1364 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3166
timestamp 1681620392
transform 1 0 1220 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3167
timestamp 1681620392
transform 1 0 1260 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3190
timestamp 1681620392
transform 1 0 1332 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3102
timestamp 1681620392
transform 1 0 1404 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3718
timestamp 1681620392
transform 1 0 1396 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3719
timestamp 1681620392
transform 1 0 1404 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_3191
timestamp 1681620392
transform 1 0 1412 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3207
timestamp 1681620392
transform 1 0 1404 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3080
timestamp 1681620392
transform 1 0 1444 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3103
timestamp 1681620392
transform 1 0 1452 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3587
timestamp 1681620392
transform 1 0 1444 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_3142
timestamp 1681620392
transform 1 0 1468 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3104
timestamp 1681620392
transform 1 0 1484 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3588
timestamp 1681620392
transform 1 0 1492 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3671
timestamp 1681620392
transform 1 0 1476 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3672
timestamp 1681620392
transform 1 0 1484 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3168
timestamp 1681620392
transform 1 0 1476 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3192
timestamp 1681620392
transform 1 0 1468 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3143
timestamp 1681620392
transform 1 0 1492 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_3673
timestamp 1681620392
transform 1 0 1500 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3081
timestamp 1681620392
transform 1 0 1540 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_3555
timestamp 1681620392
transform 1 0 1532 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_3589
timestamp 1681620392
transform 1 0 1540 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3674
timestamp 1681620392
transform 1 0 1548 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3675
timestamp 1681620392
transform 1 0 1556 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3169
timestamp 1681620392
transform 1 0 1556 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3193
timestamp 1681620392
transform 1 0 1548 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3082
timestamp 1681620392
transform 1 0 1604 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3105
timestamp 1681620392
transform 1 0 1580 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3083
timestamp 1681620392
transform 1 0 1620 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_3590
timestamp 1681620392
transform 1 0 1580 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3591
timestamp 1681620392
transform 1 0 1596 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3592
timestamp 1681620392
transform 1 0 1612 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3676
timestamp 1681620392
transform 1 0 1588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3677
timestamp 1681620392
transform 1 0 1604 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3678
timestamp 1681620392
transform 1 0 1620 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3194
timestamp 1681620392
transform 1 0 1620 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3106
timestamp 1681620392
transform 1 0 1660 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3593
timestamp 1681620392
transform 1 0 1652 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3679
timestamp 1681620392
transform 1 0 1652 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3594
timestamp 1681620392
transform 1 0 1684 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3680
timestamp 1681620392
transform 1 0 1676 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3107
timestamp 1681620392
transform 1 0 1692 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3681
timestamp 1681620392
transform 1 0 1724 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3720
timestamp 1681620392
transform 1 0 1748 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3595
timestamp 1681620392
transform 1 0 1764 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_3067
timestamp 1681620392
transform 1 0 1804 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3068
timestamp 1681620392
transform 1 0 1836 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_3596
timestamp 1681620392
transform 1 0 1780 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_3130
timestamp 1681620392
transform 1 0 1828 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_3682
timestamp 1681620392
transform 1 0 1828 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3084
timestamp 1681620392
transform 1 0 1876 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3131
timestamp 1681620392
transform 1 0 1884 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_3597
timestamp 1681620392
transform 1 0 1900 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_3144
timestamp 1681620392
transform 1 0 1892 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3170
timestamp 1681620392
transform 1 0 1900 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_3598
timestamp 1681620392
transform 1 0 1924 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_3171
timestamp 1681620392
transform 1 0 1932 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_3599
timestamp 1681620392
transform 1 0 1964 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3721
timestamp 1681620392
transform 1 0 1964 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_3208
timestamp 1681620392
transform 1 0 1964 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3108
timestamp 1681620392
transform 1 0 1996 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3600
timestamp 1681620392
transform 1 0 1996 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_3069
timestamp 1681620392
transform 1 0 2012 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3070
timestamp 1681620392
transform 1 0 2044 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3085
timestamp 1681620392
transform 1 0 2100 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3109
timestamp 1681620392
transform 1 0 2028 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3110
timestamp 1681620392
transform 1 0 2060 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3111
timestamp 1681620392
transform 1 0 2116 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3601
timestamp 1681620392
transform 1 0 2012 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3602
timestamp 1681620392
transform 1 0 2100 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3603
timestamp 1681620392
transform 1 0 2116 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3604
timestamp 1681620392
transform 1 0 2132 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3605
timestamp 1681620392
transform 1 0 2140 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3683
timestamp 1681620392
transform 1 0 2060 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3684
timestamp 1681620392
transform 1 0 2092 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3685
timestamp 1681620392
transform 1 0 2108 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3686
timestamp 1681620392
transform 1 0 2124 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3145
timestamp 1681620392
transform 1 0 2132 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3172
timestamp 1681620392
transform 1 0 2140 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3071
timestamp 1681620392
transform 1 0 2180 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3112
timestamp 1681620392
transform 1 0 2164 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3113
timestamp 1681620392
transform 1 0 2204 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3606
timestamp 1681620392
transform 1 0 2164 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3607
timestamp 1681620392
transform 1 0 2180 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3608
timestamp 1681620392
transform 1 0 2268 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3687
timestamp 1681620392
transform 1 0 2204 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3688
timestamp 1681620392
transform 1 0 2260 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3689
timestamp 1681620392
transform 1 0 2268 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3722
timestamp 1681620392
transform 1 0 2164 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_3173
timestamp 1681620392
transform 1 0 2180 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3174
timestamp 1681620392
transform 1 0 2260 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3195
timestamp 1681620392
transform 1 0 2164 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3196
timestamp 1681620392
transform 1 0 2268 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3209
timestamp 1681620392
transform 1 0 2252 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3217
timestamp 1681620392
transform 1 0 2228 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_3609
timestamp 1681620392
transform 1 0 2292 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3610
timestamp 1681620392
transform 1 0 2316 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3690
timestamp 1681620392
transform 1 0 2300 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3723
timestamp 1681620392
transform 1 0 2284 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_3146
timestamp 1681620392
transform 1 0 2308 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3114
timestamp 1681620392
transform 1 0 2340 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3072
timestamp 1681620392
transform 1 0 2444 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3115
timestamp 1681620392
transform 1 0 2436 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3611
timestamp 1681620392
transform 1 0 2420 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3612
timestamp 1681620392
transform 1 0 2436 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_3116
timestamp 1681620392
transform 1 0 2516 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3613
timestamp 1681620392
transform 1 0 2452 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3614
timestamp 1681620392
transform 1 0 2476 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3615
timestamp 1681620392
transform 1 0 2484 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3616
timestamp 1681620392
transform 1 0 2508 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3617
timestamp 1681620392
transform 1 0 2516 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3691
timestamp 1681620392
transform 1 0 2324 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3692
timestamp 1681620392
transform 1 0 2340 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3693
timestamp 1681620392
transform 1 0 2396 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3694
timestamp 1681620392
transform 1 0 2436 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3695
timestamp 1681620392
transform 1 0 2444 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3724
timestamp 1681620392
transform 1 0 2308 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_3197
timestamp 1681620392
transform 1 0 2300 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3210
timestamp 1681620392
transform 1 0 2284 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3218
timestamp 1681620392
transform 1 0 2284 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3175
timestamp 1681620392
transform 1 0 2324 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_3725
timestamp 1681620392
transform 1 0 2332 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_3211
timestamp 1681620392
transform 1 0 2308 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3212
timestamp 1681620392
transform 1 0 2332 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3147
timestamp 1681620392
transform 1 0 2452 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_3696
timestamp 1681620392
transform 1 0 2468 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3697
timestamp 1681620392
transform 1 0 2500 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3726
timestamp 1681620392
transform 1 0 2452 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_3176
timestamp 1681620392
transform 1 0 2476 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_3727
timestamp 1681620392
transform 1 0 2484 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_3177
timestamp 1681620392
transform 1 0 2500 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3086
timestamp 1681620392
transform 1 0 2548 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3087
timestamp 1681620392
transform 1 0 2604 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3117
timestamp 1681620392
transform 1 0 2580 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3118
timestamp 1681620392
transform 1 0 2628 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3119
timestamp 1681620392
transform 1 0 2660 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3618
timestamp 1681620392
transform 1 0 2540 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3619
timestamp 1681620392
transform 1 0 2556 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_3132
timestamp 1681620392
transform 1 0 2588 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_3133
timestamp 1681620392
transform 1 0 2644 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_3620
timestamp 1681620392
transform 1 0 2652 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3621
timestamp 1681620392
transform 1 0 2660 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3698
timestamp 1681620392
transform 1 0 2532 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3728
timestamp 1681620392
transform 1 0 2516 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_3198
timestamp 1681620392
transform 1 0 2516 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3148
timestamp 1681620392
transform 1 0 2540 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_3699
timestamp 1681620392
transform 1 0 2580 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3149
timestamp 1681620392
transform 1 0 2628 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_3700
timestamp 1681620392
transform 1 0 2636 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3701
timestamp 1681620392
transform 1 0 2644 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3150
timestamp 1681620392
transform 1 0 2652 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3178
timestamp 1681620392
transform 1 0 2644 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_3622
timestamp 1681620392
transform 1 0 2692 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3623
timestamp 1681620392
transform 1 0 2700 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3702
timestamp 1681620392
transform 1 0 2668 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3703
timestamp 1681620392
transform 1 0 2684 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3704
timestamp 1681620392
transform 1 0 2700 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3179
timestamp 1681620392
transform 1 0 2668 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3199
timestamp 1681620392
transform 1 0 2700 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3073
timestamp 1681620392
transform 1 0 2748 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_3624
timestamp 1681620392
transform 1 0 2748 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3625
timestamp 1681620392
transform 1 0 2756 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3705
timestamp 1681620392
transform 1 0 2724 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3706
timestamp 1681620392
transform 1 0 2740 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3151
timestamp 1681620392
transform 1 0 2748 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_3707
timestamp 1681620392
transform 1 0 2756 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3180
timestamp 1681620392
transform 1 0 2724 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3200
timestamp 1681620392
transform 1 0 2756 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3120
timestamp 1681620392
transform 1 0 2772 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3152
timestamp 1681620392
transform 1 0 2772 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3201
timestamp 1681620392
transform 1 0 2780 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3134
timestamp 1681620392
transform 1 0 2788 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_3121
timestamp 1681620392
transform 1 0 2804 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3708
timestamp 1681620392
transform 1 0 2796 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_3135
timestamp 1681620392
transform 1 0 2828 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_3202
timestamp 1681620392
transform 1 0 2820 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3213
timestamp 1681620392
transform 1 0 2836 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_3626
timestamp 1681620392
transform 1 0 2860 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_3153
timestamp 1681620392
transform 1 0 2860 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3088
timestamp 1681620392
transform 1 0 2892 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3122
timestamp 1681620392
transform 1 0 2884 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3123
timestamp 1681620392
transform 1 0 2924 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_3627
timestamp 1681620392
transform 1 0 2884 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3628
timestamp 1681620392
transform 1 0 2892 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3629
timestamp 1681620392
transform 1 0 2916 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3630
timestamp 1681620392
transform 1 0 2924 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3709
timestamp 1681620392
transform 1 0 2876 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3710
timestamp 1681620392
transform 1 0 2892 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3711
timestamp 1681620392
transform 1 0 2908 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3712
timestamp 1681620392
transform 1 0 2924 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3729
timestamp 1681620392
transform 1 0 2860 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_3181
timestamp 1681620392
transform 1 0 2868 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3182
timestamp 1681620392
transform 1 0 2892 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3203
timestamp 1681620392
transform 1 0 2924 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3214
timestamp 1681620392
transform 1 0 2924 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_3631
timestamp 1681620392
transform 1 0 2948 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_3154
timestamp 1681620392
transform 1 0 2948 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_3632
timestamp 1681620392
transform 1 0 2996 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3713
timestamp 1681620392
transform 1 0 3004 0 1 1125
box -2 -2 2 2
use Project_Top_VIA0  Project_Top_VIA0_38
timestamp 1681620392
transform 1 0 24 0 1 1070
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_194
timestamp 1681620392
transform 1 0 72 0 -1 1170
box -8 -3 104 105
use FILL  FILL_818
timestamp 1681620392
transform 1 0 168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_820
timestamp 1681620392
transform 1 0 176 0 -1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_83
timestamp 1681620392
transform 1 0 184 0 -1 1170
box -8 -3 40 105
use INVX2  INVX2_239
timestamp 1681620392
transform 1 0 216 0 -1 1170
box -9 -3 26 105
use FILL  FILL_835
timestamp 1681620392
transform 1 0 232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_836
timestamp 1681620392
transform 1 0 240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_837
timestamp 1681620392
transform 1 0 248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_838
timestamp 1681620392
transform 1 0 256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_839
timestamp 1681620392
transform 1 0 264 0 -1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_72
timestamp 1681620392
transform 1 0 272 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_73
timestamp 1681620392
transform 1 0 296 0 -1 1170
box -8 -3 32 105
use INVX2  INVX2_240
timestamp 1681620392
transform 1 0 320 0 -1 1170
box -9 -3 26 105
use FILL  FILL_840
timestamp 1681620392
transform 1 0 336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_841
timestamp 1681620392
transform 1 0 344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_842
timestamp 1681620392
transform 1 0 352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_843
timestamp 1681620392
transform 1 0 360 0 -1 1170
box -8 -3 16 105
use FILL  FILL_844
timestamp 1681620392
transform 1 0 368 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_63
timestamp 1681620392
transform -1 0 416 0 -1 1170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_208
timestamp 1681620392
transform -1 0 512 0 -1 1170
box -8 -3 104 105
use OAI22X1  OAI22X1_64
timestamp 1681620392
transform -1 0 552 0 -1 1170
box -8 -3 46 105
use OAI21X1  OAI21X1_210
timestamp 1681620392
transform -1 0 584 0 -1 1170
box -8 -3 34 105
use FILL  FILL_845
timestamp 1681620392
transform 1 0 584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_846
timestamp 1681620392
transform 1 0 592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_847
timestamp 1681620392
transform 1 0 600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_848
timestamp 1681620392
transform 1 0 608 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_241
timestamp 1681620392
transform 1 0 616 0 -1 1170
box -9 -3 26 105
use FILL  FILL_849
timestamp 1681620392
transform 1 0 632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_850
timestamp 1681620392
transform 1 0 640 0 -1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_211
timestamp 1681620392
transform -1 0 680 0 -1 1170
box -8 -3 34 105
use FILL  FILL_851
timestamp 1681620392
transform 1 0 680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_852
timestamp 1681620392
transform 1 0 688 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_242
timestamp 1681620392
transform -1 0 712 0 -1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_209
timestamp 1681620392
transform 1 0 712 0 -1 1170
box -8 -3 104 105
use FILL  FILL_853
timestamp 1681620392
transform 1 0 808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_854
timestamp 1681620392
transform 1 0 816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_855
timestamp 1681620392
transform 1 0 824 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_3219
timestamp 1681620392
transform 1 0 868 0 1 1075
box -3 -3 3 3
use AOI22X1  AOI22X1_26
timestamp 1681620392
transform 1 0 832 0 -1 1170
box -8 -3 46 105
use FILL  FILL_856
timestamp 1681620392
transform 1 0 872 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_27
timestamp 1681620392
transform -1 0 920 0 -1 1170
box -8 -3 46 105
use FILL  FILL_857
timestamp 1681620392
transform 1 0 920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_858
timestamp 1681620392
transform 1 0 928 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_3220
timestamp 1681620392
transform 1 0 1020 0 1 1075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_210
timestamp 1681620392
transform 1 0 936 0 -1 1170
box -8 -3 104 105
use INVX2  INVX2_243
timestamp 1681620392
transform 1 0 1032 0 -1 1170
box -9 -3 26 105
use AOI21X1  AOI21X1_22
timestamp 1681620392
transform -1 0 1080 0 -1 1170
box -7 -3 39 105
use DFFNEGX1  DFFNEGX1_211
timestamp 1681620392
transform 1 0 1080 0 -1 1170
box -8 -3 104 105
use FILL  FILL_859
timestamp 1681620392
transform 1 0 1176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_860
timestamp 1681620392
transform 1 0 1184 0 -1 1170
box -8 -3 16 105
use AOI21X1  AOI21X1_23
timestamp 1681620392
transform 1 0 1192 0 -1 1170
box -7 -3 39 105
use DFFNEGX1  DFFNEGX1_212
timestamp 1681620392
transform 1 0 1224 0 -1 1170
box -8 -3 104 105
use OAI22X1  OAI22X1_65
timestamp 1681620392
transform 1 0 1320 0 -1 1170
box -8 -3 46 105
use NAND2X1  NAND2X1_213
timestamp 1681620392
transform 1 0 1360 0 -1 1170
box -8 -3 32 105
use FILL  FILL_861
timestamp 1681620392
transform 1 0 1384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_862
timestamp 1681620392
transform 1 0 1392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_863
timestamp 1681620392
transform 1 0 1400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_864
timestamp 1681620392
transform 1 0 1408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_865
timestamp 1681620392
transform 1 0 1416 0 -1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_214
timestamp 1681620392
transform -1 0 1448 0 -1 1170
box -8 -3 32 105
use FILL  FILL_866
timestamp 1681620392
transform 1 0 1448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_867
timestamp 1681620392
transform 1 0 1456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_868
timestamp 1681620392
transform 1 0 1464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_869
timestamp 1681620392
transform 1 0 1472 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_244
timestamp 1681620392
transform -1 0 1496 0 -1 1170
box -9 -3 26 105
use OR2X1  OR2X1_6
timestamp 1681620392
transform -1 0 1528 0 -1 1170
box -8 -3 40 105
use FILL  FILL_870
timestamp 1681620392
transform 1 0 1528 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_245
timestamp 1681620392
transform 1 0 1536 0 -1 1170
box -9 -3 26 105
use FILL  FILL_871
timestamp 1681620392
transform 1 0 1552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_872
timestamp 1681620392
transform 1 0 1560 0 -1 1170
box -8 -3 16 105
use FILL  FILL_873
timestamp 1681620392
transform 1 0 1568 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_66
timestamp 1681620392
transform 1 0 1576 0 -1 1170
box -8 -3 46 105
use FILL  FILL_874
timestamp 1681620392
transform 1 0 1616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_875
timestamp 1681620392
transform 1 0 1624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_876
timestamp 1681620392
transform 1 0 1632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_877
timestamp 1681620392
transform 1 0 1640 0 -1 1170
box -8 -3 16 105
use AOI21X1  AOI21X1_24
timestamp 1681620392
transform 1 0 1648 0 -1 1170
box -7 -3 39 105
use INVX2  INVX2_246
timestamp 1681620392
transform 1 0 1680 0 -1 1170
box -9 -3 26 105
use FILL  FILL_878
timestamp 1681620392
transform 1 0 1696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_879
timestamp 1681620392
transform 1 0 1704 0 -1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_212
timestamp 1681620392
transform 1 0 1712 0 -1 1170
box -8 -3 34 105
use FILL  FILL_880
timestamp 1681620392
transform 1 0 1744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_881
timestamp 1681620392
transform 1 0 1752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_882
timestamp 1681620392
transform 1 0 1760 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_213
timestamp 1681620392
transform 1 0 1768 0 -1 1170
box -8 -3 104 105
use INVX2  INVX2_247
timestamp 1681620392
transform 1 0 1864 0 -1 1170
box -9 -3 26 105
use FILL  FILL_883
timestamp 1681620392
transform 1 0 1880 0 -1 1170
box -8 -3 16 105
use FILL  FILL_884
timestamp 1681620392
transform 1 0 1888 0 -1 1170
box -8 -3 16 105
use FILL  FILL_885
timestamp 1681620392
transform 1 0 1896 0 -1 1170
box -8 -3 16 105
use FILL  FILL_886
timestamp 1681620392
transform 1 0 1904 0 -1 1170
box -8 -3 16 105
use FILL  FILL_887
timestamp 1681620392
transform 1 0 1912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_888
timestamp 1681620392
transform 1 0 1920 0 -1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_213
timestamp 1681620392
transform 1 0 1928 0 -1 1170
box -8 -3 34 105
use NAND2X1  NAND2X1_215
timestamp 1681620392
transform -1 0 1984 0 -1 1170
box -8 -3 32 105
use FILL  FILL_889
timestamp 1681620392
transform 1 0 1984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_890
timestamp 1681620392
transform 1 0 1992 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_214
timestamp 1681620392
transform 1 0 2000 0 -1 1170
box -8 -3 104 105
use OAI22X1  OAI22X1_67
timestamp 1681620392
transform -1 0 2136 0 -1 1170
box -8 -3 46 105
use OAI21X1  OAI21X1_214
timestamp 1681620392
transform 1 0 2136 0 -1 1170
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_215
timestamp 1681620392
transform 1 0 2168 0 -1 1170
box -8 -3 104 105
use NAND2X1  NAND2X1_216
timestamp 1681620392
transform 1 0 2264 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_217
timestamp 1681620392
transform 1 0 2288 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_218
timestamp 1681620392
transform 1 0 2312 0 -1 1170
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_216
timestamp 1681620392
transform -1 0 2432 0 -1 1170
box -8 -3 104 105
use INVX2  INVX2_248
timestamp 1681620392
transform 1 0 2432 0 -1 1170
box -9 -3 26 105
use OAI21X1  OAI21X1_215
timestamp 1681620392
transform -1 0 2480 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_216
timestamp 1681620392
transform -1 0 2512 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_217
timestamp 1681620392
transform -1 0 2544 0 -1 1170
box -8 -3 34 105
use M3_M2  M3_M2_3221
timestamp 1681620392
transform 1 0 2604 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3222
timestamp 1681620392
transform 1 0 2620 0 1 1075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_217
timestamp 1681620392
transform 1 0 2544 0 -1 1170
box -8 -3 104 105
use INVX2  INVX2_249
timestamp 1681620392
transform -1 0 2656 0 -1 1170
box -9 -3 26 105
use FILL  FILL_891
timestamp 1681620392
transform 1 0 2656 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_28
timestamp 1681620392
transform -1 0 2704 0 -1 1170
box -8 -3 46 105
use FILL  FILL_892
timestamp 1681620392
transform 1 0 2704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_898
timestamp 1681620392
transform 1 0 2712 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_30
timestamp 1681620392
transform -1 0 2760 0 -1 1170
box -8 -3 46 105
use FILL  FILL_899
timestamp 1681620392
transform 1 0 2760 0 -1 1170
box -8 -3 16 105
use FILL  FILL_900
timestamp 1681620392
transform 1 0 2768 0 -1 1170
box -8 -3 16 105
use FILL  FILL_901
timestamp 1681620392
transform 1 0 2776 0 -1 1170
box -8 -3 16 105
use FILL  FILL_902
timestamp 1681620392
transform 1 0 2784 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_250
timestamp 1681620392
transform 1 0 2792 0 -1 1170
box -9 -3 26 105
use FILL  FILL_903
timestamp 1681620392
transform 1 0 2808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_904
timestamp 1681620392
transform 1 0 2816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_905
timestamp 1681620392
transform 1 0 2824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_906
timestamp 1681620392
transform 1 0 2832 0 -1 1170
box -8 -3 16 105
use FILL  FILL_907
timestamp 1681620392
transform 1 0 2840 0 -1 1170
box -8 -3 16 105
use FILL  FILL_908
timestamp 1681620392
transform 1 0 2848 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_3223
timestamp 1681620392
transform 1 0 2868 0 1 1075
box -3 -3 3 3
use OAI21X1  OAI21X1_220
timestamp 1681620392
transform -1 0 2888 0 -1 1170
box -8 -3 34 105
use AOI22X1  AOI22X1_31
timestamp 1681620392
transform 1 0 2888 0 -1 1170
box -8 -3 46 105
use INVX2  INVX2_251
timestamp 1681620392
transform 1 0 2928 0 -1 1170
box -9 -3 26 105
use FILL  FILL_909
timestamp 1681620392
transform 1 0 2944 0 -1 1170
box -8 -3 16 105
use FILL  FILL_910
timestamp 1681620392
transform 1 0 2952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_917
timestamp 1681620392
transform 1 0 2960 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_3224
timestamp 1681620392
transform 1 0 2980 0 1 1075
box -3 -3 3 3
use OAI21X1  OAI21X1_221
timestamp 1681620392
transform -1 0 3000 0 -1 1170
box -8 -3 34 105
use FILL  FILL_918
timestamp 1681620392
transform 1 0 3000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_920
timestamp 1681620392
transform 1 0 3008 0 -1 1170
box -8 -3 16 105
use Project_Top_VIA0  Project_Top_VIA0_39
timestamp 1681620392
transform 1 0 3067 0 1 1070
box -10 -3 10 3
use M3_M2  M3_M2_3333
timestamp 1681620392
transform 1 0 68 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3308
timestamp 1681620392
transform 1 0 124 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3250
timestamp 1681620392
transform 1 0 164 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3275
timestamp 1681620392
transform 1 0 140 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3761
timestamp 1681620392
transform 1 0 140 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3762
timestamp 1681620392
transform 1 0 156 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3309
timestamp 1681620392
transform 1 0 164 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_3763
timestamp 1681620392
transform 1 0 172 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3850
timestamp 1681620392
transform 1 0 132 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3851
timestamp 1681620392
transform 1 0 148 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3334
timestamp 1681620392
transform 1 0 156 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_3852
timestamp 1681620392
transform 1 0 164 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3380
timestamp 1681620392
transform 1 0 132 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3351
timestamp 1681620392
transform 1 0 164 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3276
timestamp 1681620392
transform 1 0 180 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3853
timestamp 1681620392
transform 1 0 180 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3854
timestamp 1681620392
transform 1 0 188 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3352
timestamp 1681620392
transform 1 0 188 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3251
timestamp 1681620392
transform 1 0 204 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3277
timestamp 1681620392
transform 1 0 212 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3764
timestamp 1681620392
transform 1 0 212 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3932
timestamp 1681620392
transform 1 0 236 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_3381
timestamp 1681620392
transform 1 0 236 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3278
timestamp 1681620392
transform 1 0 252 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3765
timestamp 1681620392
transform 1 0 252 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3239
timestamp 1681620392
transform 1 0 292 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_3766
timestamp 1681620392
transform 1 0 284 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3855
timestamp 1681620392
transform 1 0 260 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3856
timestamp 1681620392
transform 1 0 268 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3857
timestamp 1681620392
transform 1 0 276 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3933
timestamp 1681620392
transform 1 0 252 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_3382
timestamp 1681620392
transform 1 0 252 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3383
timestamp 1681620392
transform 1 0 268 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3353
timestamp 1681620392
transform 1 0 284 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_3767
timestamp 1681620392
transform 1 0 308 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3279
timestamp 1681620392
transform 1 0 340 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3734
timestamp 1681620392
transform 1 0 348 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3768
timestamp 1681620392
transform 1 0 340 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3858
timestamp 1681620392
transform 1 0 316 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3859
timestamp 1681620392
transform 1 0 324 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3354
timestamp 1681620392
transform 1 0 316 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_3934
timestamp 1681620392
transform 1 0 340 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_3384
timestamp 1681620392
transform 1 0 324 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3240
timestamp 1681620392
transform 1 0 380 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3252
timestamp 1681620392
transform 1 0 372 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_3769
timestamp 1681620392
transform 1 0 372 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3860
timestamp 1681620392
transform 1 0 364 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3355
timestamp 1681620392
transform 1 0 364 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3385
timestamp 1681620392
transform 1 0 356 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_3735
timestamp 1681620392
transform 1 0 388 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3770
timestamp 1681620392
transform 1 0 388 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3335
timestamp 1681620392
transform 1 0 388 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_3861
timestamp 1681620392
transform 1 0 396 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3356
timestamp 1681620392
transform 1 0 396 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3253
timestamp 1681620392
transform 1 0 420 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_3731
timestamp 1681620392
transform 1 0 428 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_3736
timestamp 1681620392
transform 1 0 412 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3737
timestamp 1681620392
transform 1 0 420 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_3280
timestamp 1681620392
transform 1 0 428 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3254
timestamp 1681620392
transform 1 0 460 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_3732
timestamp 1681620392
transform 1 0 484 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_3738
timestamp 1681620392
transform 1 0 452 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3771
timestamp 1681620392
transform 1 0 412 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3310
timestamp 1681620392
transform 1 0 420 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_3772
timestamp 1681620392
transform 1 0 428 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3386
timestamp 1681620392
transform 1 0 404 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_3739
timestamp 1681620392
transform 1 0 484 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3773
timestamp 1681620392
transform 1 0 460 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3774
timestamp 1681620392
transform 1 0 476 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3862
timestamp 1681620392
transform 1 0 452 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3387
timestamp 1681620392
transform 1 0 436 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3311
timestamp 1681620392
transform 1 0 484 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3255
timestamp 1681620392
transform 1 0 532 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3256
timestamp 1681620392
transform 1 0 564 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_3740
timestamp 1681620392
transform 1 0 508 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3775
timestamp 1681620392
transform 1 0 492 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3336
timestamp 1681620392
transform 1 0 492 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_3776
timestamp 1681620392
transform 1 0 524 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3777
timestamp 1681620392
transform 1 0 564 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3312
timestamp 1681620392
transform 1 0 580 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3281
timestamp 1681620392
transform 1 0 668 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3778
timestamp 1681620392
transform 1 0 620 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3779
timestamp 1681620392
transform 1 0 660 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3780
timestamp 1681620392
transform 1 0 716 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3781
timestamp 1681620392
transform 1 0 724 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3782
timestamp 1681620392
transform 1 0 732 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3783
timestamp 1681620392
transform 1 0 740 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3863
timestamp 1681620392
transform 1 0 516 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3337
timestamp 1681620392
transform 1 0 524 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_3864
timestamp 1681620392
transform 1 0 540 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3357
timestamp 1681620392
transform 1 0 540 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_3865
timestamp 1681620392
transform 1 0 636 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3866
timestamp 1681620392
transform 1 0 724 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3358
timestamp 1681620392
transform 1 0 636 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3282
timestamp 1681620392
transform 1 0 764 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3784
timestamp 1681620392
transform 1 0 764 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3867
timestamp 1681620392
transform 1 0 764 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3359
timestamp 1681620392
transform 1 0 764 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_3785
timestamp 1681620392
transform 1 0 812 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3868
timestamp 1681620392
transform 1 0 804 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3257
timestamp 1681620392
transform 1 0 844 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_3786
timestamp 1681620392
transform 1 0 828 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3787
timestamp 1681620392
transform 1 0 844 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3869
timestamp 1681620392
transform 1 0 820 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3388
timestamp 1681620392
transform 1 0 812 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3313
timestamp 1681620392
transform 1 0 852 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3225
timestamp 1681620392
transform 1 0 932 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_3230
timestamp 1681620392
transform 1 0 924 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3241
timestamp 1681620392
transform 1 0 900 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3258
timestamp 1681620392
transform 1 0 892 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3283
timestamp 1681620392
transform 1 0 876 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3741
timestamp 1681620392
transform 1 0 892 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_3284
timestamp 1681620392
transform 1 0 940 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3788
timestamp 1681620392
transform 1 0 868 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3789
timestamp 1681620392
transform 1 0 876 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3790
timestamp 1681620392
transform 1 0 892 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3791
timestamp 1681620392
transform 1 0 916 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3792
timestamp 1681620392
transform 1 0 932 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3793
timestamp 1681620392
transform 1 0 940 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3338
timestamp 1681620392
transform 1 0 844 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_3870
timestamp 1681620392
transform 1 0 852 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3871
timestamp 1681620392
transform 1 0 860 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3872
timestamp 1681620392
transform 1 0 892 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3339
timestamp 1681620392
transform 1 0 900 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_3873
timestamp 1681620392
transform 1 0 908 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3874
timestamp 1681620392
transform 1 0 924 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3875
timestamp 1681620392
transform 1 0 932 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3360
timestamp 1681620392
transform 1 0 860 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3361
timestamp 1681620392
transform 1 0 876 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3362
timestamp 1681620392
transform 1 0 892 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3231
timestamp 1681620392
transform 1 0 980 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3242
timestamp 1681620392
transform 1 0 980 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_3742
timestamp 1681620392
transform 1 0 980 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_3314
timestamp 1681620392
transform 1 0 988 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_3876
timestamp 1681620392
transform 1 0 980 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3363
timestamp 1681620392
transform 1 0 980 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_3877
timestamp 1681620392
transform 1 0 988 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3389
timestamp 1681620392
transform 1 0 988 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3340
timestamp 1681620392
transform 1 0 1004 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3390
timestamp 1681620392
transform 1 0 1004 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3226
timestamp 1681620392
transform 1 0 1052 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_3243
timestamp 1681620392
transform 1 0 1052 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3259
timestamp 1681620392
transform 1 0 1036 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3285
timestamp 1681620392
transform 1 0 1060 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3794
timestamp 1681620392
transform 1 0 1020 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3795
timestamp 1681620392
transform 1 0 1036 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3796
timestamp 1681620392
transform 1 0 1052 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3797
timestamp 1681620392
transform 1 0 1060 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3341
timestamp 1681620392
transform 1 0 1020 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_3878
timestamp 1681620392
transform 1 0 1044 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3244
timestamp 1681620392
transform 1 0 1084 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3260
timestamp 1681620392
transform 1 0 1100 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_3743
timestamp 1681620392
transform 1 0 1100 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_3245
timestamp 1681620392
transform 1 0 1140 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_3798
timestamp 1681620392
transform 1 0 1100 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3799
timestamp 1681620392
transform 1 0 1124 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3800
timestamp 1681620392
transform 1 0 1140 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3801
timestamp 1681620392
transform 1 0 1156 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3879
timestamp 1681620392
transform 1 0 1076 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3342
timestamp 1681620392
transform 1 0 1100 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_3880
timestamp 1681620392
transform 1 0 1108 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3881
timestamp 1681620392
transform 1 0 1116 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3882
timestamp 1681620392
transform 1 0 1140 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3286
timestamp 1681620392
transform 1 0 1204 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3287
timestamp 1681620392
transform 1 0 1268 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3802
timestamp 1681620392
transform 1 0 1172 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3883
timestamp 1681620392
transform 1 0 1164 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3315
timestamp 1681620392
transform 1 0 1204 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_3803
timestamp 1681620392
transform 1 0 1228 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3316
timestamp 1681620392
transform 1 0 1252 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_3804
timestamp 1681620392
transform 1 0 1268 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3884
timestamp 1681620392
transform 1 0 1252 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3288
timestamp 1681620392
transform 1 0 1292 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3289
timestamp 1681620392
transform 1 0 1316 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3805
timestamp 1681620392
transform 1 0 1300 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3806
timestamp 1681620392
transform 1 0 1316 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3885
timestamp 1681620392
transform 1 0 1292 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3290
timestamp 1681620392
transform 1 0 1340 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3317
timestamp 1681620392
transform 1 0 1340 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_3886
timestamp 1681620392
transform 1 0 1308 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3887
timestamp 1681620392
transform 1 0 1324 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3888
timestamp 1681620392
transform 1 0 1332 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3391
timestamp 1681620392
transform 1 0 1324 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3291
timestamp 1681620392
transform 1 0 1388 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3318
timestamp 1681620392
transform 1 0 1364 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_3807
timestamp 1681620392
transform 1 0 1388 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3319
timestamp 1681620392
transform 1 0 1428 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_3889
timestamp 1681620392
transform 1 0 1364 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3292
timestamp 1681620392
transform 1 0 1476 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3808
timestamp 1681620392
transform 1 0 1468 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3293
timestamp 1681620392
transform 1 0 1500 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3809
timestamp 1681620392
transform 1 0 1484 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3810
timestamp 1681620392
transform 1 0 1500 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3811
timestamp 1681620392
transform 1 0 1524 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3890
timestamp 1681620392
transform 1 0 1492 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3891
timestamp 1681620392
transform 1 0 1508 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3892
timestamp 1681620392
transform 1 0 1516 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3364
timestamp 1681620392
transform 1 0 1508 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_3812
timestamp 1681620392
transform 1 0 1548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3935
timestamp 1681620392
transform 1 0 1564 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_3227
timestamp 1681620392
transform 1 0 1596 0 1 1065
box -3 -3 3 3
use M2_M1  M2_M1_3744
timestamp 1681620392
transform 1 0 1588 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_3320
timestamp 1681620392
transform 1 0 1588 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3294
timestamp 1681620392
transform 1 0 1612 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3813
timestamp 1681620392
transform 1 0 1604 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3893
timestamp 1681620392
transform 1 0 1588 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3894
timestamp 1681620392
transform 1 0 1612 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3246
timestamp 1681620392
transform 1 0 1636 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3232
timestamp 1681620392
transform 1 0 1652 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_3895
timestamp 1681620392
transform 1 0 1644 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3365
timestamp 1681620392
transform 1 0 1644 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3261
timestamp 1681620392
transform 1 0 1676 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_3745
timestamp 1681620392
transform 1 0 1676 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3814
timestamp 1681620392
transform 1 0 1660 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3247
timestamp 1681620392
transform 1 0 1692 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_3746
timestamp 1681620392
transform 1 0 1692 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_3321
timestamp 1681620392
transform 1 0 1684 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3233
timestamp 1681620392
transform 1 0 1724 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3262
timestamp 1681620392
transform 1 0 1716 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3263
timestamp 1681620392
transform 1 0 1732 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_3733
timestamp 1681620392
transform 1 0 1740 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_3747
timestamp 1681620392
transform 1 0 1716 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3748
timestamp 1681620392
transform 1 0 1724 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3815
timestamp 1681620392
transform 1 0 1692 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3816
timestamp 1681620392
transform 1 0 1708 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3896
timestamp 1681620392
transform 1 0 1668 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3343
timestamp 1681620392
transform 1 0 1684 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3344
timestamp 1681620392
transform 1 0 1700 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3366
timestamp 1681620392
transform 1 0 1668 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3367
timestamp 1681620392
transform 1 0 1692 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3295
timestamp 1681620392
transform 1 0 1740 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3749
timestamp 1681620392
transform 1 0 1748 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3897
timestamp 1681620392
transform 1 0 1732 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3368
timestamp 1681620392
transform 1 0 1724 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3234
timestamp 1681620392
transform 1 0 1868 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_3817
timestamp 1681620392
transform 1 0 1812 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3818
timestamp 1681620392
transform 1 0 1860 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3819
timestamp 1681620392
transform 1 0 1868 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3898
timestamp 1681620392
transform 1 0 1780 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3899
timestamp 1681620392
transform 1 0 1868 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3369
timestamp 1681620392
transform 1 0 1780 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_3750
timestamp 1681620392
transform 1 0 1908 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3820
timestamp 1681620392
transform 1 0 1900 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3322
timestamp 1681620392
transform 1 0 1908 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3345
timestamp 1681620392
transform 1 0 1900 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3264
timestamp 1681620392
transform 1 0 1924 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3265
timestamp 1681620392
transform 1 0 2004 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3296
timestamp 1681620392
transform 1 0 1924 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3297
timestamp 1681620392
transform 1 0 1956 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3821
timestamp 1681620392
transform 1 0 1972 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3323
timestamp 1681620392
transform 1 0 1988 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_3900
timestamp 1681620392
transform 1 0 1924 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3370
timestamp 1681620392
transform 1 0 1924 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3371
timestamp 1681620392
transform 1 0 1948 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3372
timestamp 1681620392
transform 1 0 1972 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3228
timestamp 1681620392
transform 1 0 2020 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_3298
timestamp 1681620392
transform 1 0 2028 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3299
timestamp 1681620392
transform 1 0 2044 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3324
timestamp 1681620392
transform 1 0 2036 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_3822
timestamp 1681620392
transform 1 0 2044 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3823
timestamp 1681620392
transform 1 0 2060 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3325
timestamp 1681620392
transform 1 0 2068 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_3901
timestamp 1681620392
transform 1 0 2036 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3902
timestamp 1681620392
transform 1 0 2052 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3346
timestamp 1681620392
transform 1 0 2060 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_3903
timestamp 1681620392
transform 1 0 2068 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3373
timestamp 1681620392
transform 1 0 2052 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3392
timestamp 1681620392
transform 1 0 2028 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3326
timestamp 1681620392
transform 1 0 2084 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_3824
timestamp 1681620392
transform 1 0 2092 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3229
timestamp 1681620392
transform 1 0 2108 0 1 1065
box -3 -3 3 3
use M2_M1  M2_M1_3904
timestamp 1681620392
transform 1 0 2100 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3825
timestamp 1681620392
transform 1 0 2124 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3905
timestamp 1681620392
transform 1 0 2124 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3300
timestamp 1681620392
transform 1 0 2148 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3826
timestamp 1681620392
transform 1 0 2140 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3827
timestamp 1681620392
transform 1 0 2148 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3235
timestamp 1681620392
transform 1 0 2172 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_3906
timestamp 1681620392
transform 1 0 2156 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3907
timestamp 1681620392
transform 1 0 2164 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3236
timestamp 1681620392
transform 1 0 2220 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3266
timestamp 1681620392
transform 1 0 2196 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_3751
timestamp 1681620392
transform 1 0 2196 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_3267
timestamp 1681620392
transform 1 0 2308 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_3752
timestamp 1681620392
transform 1 0 2300 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3828
timestamp 1681620392
transform 1 0 2236 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3829
timestamp 1681620392
transform 1 0 2300 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3830
timestamp 1681620392
transform 1 0 2308 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3908
timestamp 1681620392
transform 1 0 2196 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3909
timestamp 1681620392
transform 1 0 2212 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3374
timestamp 1681620392
transform 1 0 2196 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3375
timestamp 1681620392
transform 1 0 2236 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3393
timestamp 1681620392
transform 1 0 2212 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_3910
timestamp 1681620392
transform 1 0 2316 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3911
timestamp 1681620392
transform 1 0 2324 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3237
timestamp 1681620392
transform 1 0 2348 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3268
timestamp 1681620392
transform 1 0 2340 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_3753
timestamp 1681620392
transform 1 0 2340 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3831
timestamp 1681620392
transform 1 0 2348 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3912
timestamp 1681620392
transform 1 0 2340 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3269
timestamp 1681620392
transform 1 0 2364 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_3754
timestamp 1681620392
transform 1 0 2364 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3913
timestamp 1681620392
transform 1 0 2396 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3327
timestamp 1681620392
transform 1 0 2420 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_3914
timestamp 1681620392
transform 1 0 2436 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3832
timestamp 1681620392
transform 1 0 2460 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3238
timestamp 1681620392
transform 1 0 2484 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3301
timestamp 1681620392
transform 1 0 2508 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3328
timestamp 1681620392
transform 1 0 2476 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3302
timestamp 1681620392
transform 1 0 2564 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3833
timestamp 1681620392
transform 1 0 2500 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3834
timestamp 1681620392
transform 1 0 2556 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3835
timestamp 1681620392
transform 1 0 2564 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3915
timestamp 1681620392
transform 1 0 2476 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3916
timestamp 1681620392
transform 1 0 2572 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3376
timestamp 1681620392
transform 1 0 2572 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3248
timestamp 1681620392
transform 1 0 2628 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3303
timestamp 1681620392
transform 1 0 2604 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3836
timestamp 1681620392
transform 1 0 2604 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3837
timestamp 1681620392
transform 1 0 2644 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3917
timestamp 1681620392
transform 1 0 2596 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3918
timestamp 1681620392
transform 1 0 2612 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3919
timestamp 1681620392
transform 1 0 2628 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3920
timestamp 1681620392
transform 1 0 2636 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3394
timestamp 1681620392
transform 1 0 2596 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3270
timestamp 1681620392
transform 1 0 2676 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3304
timestamp 1681620392
transform 1 0 2668 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3755
timestamp 1681620392
transform 1 0 2676 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3838
timestamp 1681620392
transform 1 0 2660 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3329
timestamp 1681620392
transform 1 0 2668 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3249
timestamp 1681620392
transform 1 0 2708 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3271
timestamp 1681620392
transform 1 0 2692 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_3839
timestamp 1681620392
transform 1 0 2676 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3840
timestamp 1681620392
transform 1 0 2684 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3347
timestamp 1681620392
transform 1 0 2684 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3395
timestamp 1681620392
transform 1 0 2668 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3272
timestamp 1681620392
transform 1 0 2716 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3273
timestamp 1681620392
transform 1 0 2764 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3274
timestamp 1681620392
transform 1 0 2788 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_3756
timestamp 1681620392
transform 1 0 2732 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_3305
timestamp 1681620392
transform 1 0 2756 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3757
timestamp 1681620392
transform 1 0 2764 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3841
timestamp 1681620392
transform 1 0 2708 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3842
timestamp 1681620392
transform 1 0 2716 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3843
timestamp 1681620392
transform 1 0 2732 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3921
timestamp 1681620392
transform 1 0 2700 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3377
timestamp 1681620392
transform 1 0 2700 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3330
timestamp 1681620392
transform 1 0 2740 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3348
timestamp 1681620392
transform 1 0 2716 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_3758
timestamp 1681620392
transform 1 0 2796 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_3306
timestamp 1681620392
transform 1 0 2804 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3844
timestamp 1681620392
transform 1 0 2772 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3845
timestamp 1681620392
transform 1 0 2780 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3922
timestamp 1681620392
transform 1 0 2732 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3923
timestamp 1681620392
transform 1 0 2740 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3924
timestamp 1681620392
transform 1 0 2764 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3378
timestamp 1681620392
transform 1 0 2732 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3349
timestamp 1681620392
transform 1 0 2780 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_3925
timestamp 1681620392
transform 1 0 2796 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3396
timestamp 1681620392
transform 1 0 2796 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3331
timestamp 1681620392
transform 1 0 2812 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_3926
timestamp 1681620392
transform 1 0 2836 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3307
timestamp 1681620392
transform 1 0 2852 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_3846
timestamp 1681620392
transform 1 0 2852 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3927
timestamp 1681620392
transform 1 0 2852 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3397
timestamp 1681620392
transform 1 0 2844 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_3847
timestamp 1681620392
transform 1 0 2868 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_3332
timestamp 1681620392
transform 1 0 2876 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3350
timestamp 1681620392
transform 1 0 2876 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_3928
timestamp 1681620392
transform 1 0 2884 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3759
timestamp 1681620392
transform 1 0 2892 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3848
timestamp 1681620392
transform 1 0 2908 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3929
timestamp 1681620392
transform 1 0 2916 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_3379
timestamp 1681620392
transform 1 0 2908 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3398
timestamp 1681620392
transform 1 0 2916 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_3930
timestamp 1681620392
transform 1 0 2940 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3760
timestamp 1681620392
transform 1 0 2948 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_3399
timestamp 1681620392
transform 1 0 2948 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_3931
timestamp 1681620392
transform 1 0 2972 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3849
timestamp 1681620392
transform 1 0 2996 0 1 1015
box -2 -2 2 2
use Project_Top_VIA0  Project_Top_VIA0_40
timestamp 1681620392
transform 1 0 48 0 1 970
box -10 -3 10 3
use FILL  FILL_921
timestamp 1681620392
transform 1 0 72 0 1 970
box -8 -3 16 105
use FILL  FILL_922
timestamp 1681620392
transform 1 0 80 0 1 970
box -8 -3 16 105
use FILL  FILL_923
timestamp 1681620392
transform 1 0 88 0 1 970
box -8 -3 16 105
use FILL  FILL_924
timestamp 1681620392
transform 1 0 96 0 1 970
box -8 -3 16 105
use FILL  FILL_925
timestamp 1681620392
transform 1 0 104 0 1 970
box -8 -3 16 105
use FILL  FILL_926
timestamp 1681620392
transform 1 0 112 0 1 970
box -8 -3 16 105
use FILL  FILL_927
timestamp 1681620392
transform 1 0 120 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_70
timestamp 1681620392
transform 1 0 128 0 1 970
box -8 -3 46 105
use M3_M2  M3_M2_3400
timestamp 1681620392
transform 1 0 180 0 1 975
box -3 -3 3 3
use INVX2  INVX2_252
timestamp 1681620392
transform -1 0 184 0 1 970
box -9 -3 26 105
use FILL  FILL_928
timestamp 1681620392
transform 1 0 184 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_3401
timestamp 1681620392
transform 1 0 204 0 1 975
box -3 -3 3 3
use FILL  FILL_929
timestamp 1681620392
transform 1 0 192 0 1 970
box -8 -3 16 105
use FILL  FILL_930
timestamp 1681620392
transform 1 0 200 0 1 970
box -8 -3 16 105
use FILL  FILL_931
timestamp 1681620392
transform 1 0 208 0 1 970
box -8 -3 16 105
use INVX2  INVX2_253
timestamp 1681620392
transform 1 0 216 0 1 970
box -9 -3 26 105
use M3_M2  M3_M2_3402
timestamp 1681620392
transform 1 0 260 0 1 975
box -3 -3 3 3
use NOR2X1  NOR2X1_75
timestamp 1681620392
transform 1 0 232 0 1 970
box -8 -3 32 105
use M3_M2  M3_M2_3403
timestamp 1681620392
transform 1 0 284 0 1 975
box -3 -3 3 3
use NOR2X1  NOR2X1_77
timestamp 1681620392
transform 1 0 256 0 1 970
box -8 -3 32 105
use FILL  FILL_935
timestamp 1681620392
transform 1 0 280 0 1 970
box -8 -3 16 105
use FILL  FILL_936
timestamp 1681620392
transform 1 0 288 0 1 970
box -8 -3 16 105
use FILL  FILL_937
timestamp 1681620392
transform 1 0 296 0 1 970
box -8 -3 16 105
use FILL  FILL_938
timestamp 1681620392
transform 1 0 304 0 1 970
box -8 -3 16 105
use AOI21X1  AOI21X1_25
timestamp 1681620392
transform 1 0 312 0 1 970
box -7 -3 39 105
use M3_M2  M3_M2_3404
timestamp 1681620392
transform 1 0 372 0 1 975
box -3 -3 3 3
use NAND2X1  NAND2X1_220
timestamp 1681620392
transform -1 0 368 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_221
timestamp 1681620392
transform 1 0 368 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_222
timestamp 1681620392
transform 1 0 392 0 1 970
box -8 -3 32 105
use NAND3X1  NAND3X1_84
timestamp 1681620392
transform 1 0 416 0 1 970
box -8 -3 40 105
use AND2X2  AND2X2_22
timestamp 1681620392
transform 1 0 448 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_86
timestamp 1681620392
transform 1 0 480 0 1 970
box -8 -3 40 105
use INVX2  INVX2_255
timestamp 1681620392
transform 1 0 512 0 1 970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_219
timestamp 1681620392
transform 1 0 528 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_220
timestamp 1681620392
transform 1 0 624 0 1 970
box -8 -3 104 105
use INVX2  INVX2_256
timestamp 1681620392
transform 1 0 720 0 1 970
box -9 -3 26 105
use FILL  FILL_946
timestamp 1681620392
transform 1 0 736 0 1 970
box -8 -3 16 105
use FILL  FILL_947
timestamp 1681620392
transform 1 0 744 0 1 970
box -8 -3 16 105
use INVX2  INVX2_257
timestamp 1681620392
transform -1 0 768 0 1 970
box -9 -3 26 105
use INVX2  INVX2_258
timestamp 1681620392
transform -1 0 784 0 1 970
box -9 -3 26 105
use FILL  FILL_948
timestamp 1681620392
transform 1 0 784 0 1 970
box -8 -3 16 105
use FILL  FILL_949
timestamp 1681620392
transform 1 0 792 0 1 970
box -8 -3 16 105
use FILL  FILL_950
timestamp 1681620392
transform 1 0 800 0 1 970
box -8 -3 16 105
use FILL  FILL_951
timestamp 1681620392
transform 1 0 808 0 1 970
box -8 -3 16 105
use FILL  FILL_952
timestamp 1681620392
transform 1 0 816 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_32
timestamp 1681620392
transform 1 0 824 0 1 970
box -8 -3 46 105
use OAI21X1  OAI21X1_222
timestamp 1681620392
transform 1 0 864 0 1 970
box -8 -3 34 105
use M3_M2  M3_M2_3405
timestamp 1681620392
transform 1 0 908 0 1 975
box -3 -3 3 3
use AOI22X1  AOI22X1_33
timestamp 1681620392
transform -1 0 936 0 1 970
box -8 -3 46 105
use FILL  FILL_953
timestamp 1681620392
transform 1 0 936 0 1 970
box -8 -3 16 105
use FILL  FILL_954
timestamp 1681620392
transform 1 0 944 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_223
timestamp 1681620392
transform 1 0 952 0 1 970
box -8 -3 34 105
use FILL  FILL_955
timestamp 1681620392
transform 1 0 984 0 1 970
box -8 -3 16 105
use FILL  FILL_956
timestamp 1681620392
transform 1 0 992 0 1 970
box -8 -3 16 105
use FILL  FILL_957
timestamp 1681620392
transform 1 0 1000 0 1 970
box -8 -3 16 105
use FILL  FILL_958
timestamp 1681620392
transform 1 0 1008 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_34
timestamp 1681620392
transform -1 0 1056 0 1 970
box -8 -3 46 105
use FILL  FILL_959
timestamp 1681620392
transform 1 0 1056 0 1 970
box -8 -3 16 105
use FILL  FILL_960
timestamp 1681620392
transform 1 0 1064 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_224
timestamp 1681620392
transform 1 0 1072 0 1 970
box -8 -3 34 105
use AOI22X1  AOI22X1_35
timestamp 1681620392
transform -1 0 1144 0 1 970
box -8 -3 46 105
use INVX2  INVX2_259
timestamp 1681620392
transform -1 0 1160 0 1 970
box -9 -3 26 105
use FILL  FILL_961
timestamp 1681620392
transform 1 0 1160 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_221
timestamp 1681620392
transform -1 0 1264 0 1 970
box -8 -3 104 105
use INVX2  INVX2_260
timestamp 1681620392
transform -1 0 1280 0 1 970
box -9 -3 26 105
use FILL  FILL_962
timestamp 1681620392
transform 1 0 1280 0 1 970
box -8 -3 16 105
use FILL  FILL_974
timestamp 1681620392
transform 1 0 1288 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_36
timestamp 1681620392
transform 1 0 1296 0 1 970
box -8 -3 46 105
use FILL  FILL_976
timestamp 1681620392
transform 1 0 1336 0 1 970
box -8 -3 16 105
use FILL  FILL_978
timestamp 1681620392
transform 1 0 1344 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_224
timestamp 1681620392
transform 1 0 1352 0 1 970
box -8 -3 104 105
use FILL  FILL_979
timestamp 1681620392
transform 1 0 1448 0 1 970
box -8 -3 16 105
use INVX2  INVX2_266
timestamp 1681620392
transform 1 0 1456 0 1 970
box -9 -3 26 105
use FILL  FILL_980
timestamp 1681620392
transform 1 0 1472 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_3406
timestamp 1681620392
transform 1 0 1508 0 1 975
box -3 -3 3 3
use AOI22X1  AOI22X1_40
timestamp 1681620392
transform 1 0 1480 0 1 970
box -8 -3 46 105
use FILL  FILL_986
timestamp 1681620392
transform 1 0 1520 0 1 970
box -8 -3 16 105
use FILL  FILL_988
timestamp 1681620392
transform 1 0 1528 0 1 970
box -8 -3 16 105
use FILL  FILL_990
timestamp 1681620392
transform 1 0 1536 0 1 970
box -8 -3 16 105
use NOR2X1  NOR2X1_78
timestamp 1681620392
transform -1 0 1568 0 1 970
box -8 -3 32 105
use FILL  FILL_991
timestamp 1681620392
transform 1 0 1568 0 1 970
box -8 -3 16 105
use FILL  FILL_992
timestamp 1681620392
transform 1 0 1576 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_231
timestamp 1681620392
transform -1 0 1616 0 1 970
box -8 -3 34 105
use FILL  FILL_993
timestamp 1681620392
transform 1 0 1616 0 1 970
box -8 -3 16 105
use FILL  FILL_994
timestamp 1681620392
transform 1 0 1624 0 1 970
box -8 -3 16 105
use FILL  FILL_995
timestamp 1681620392
transform 1 0 1632 0 1 970
box -8 -3 16 105
use FILL  FILL_998
timestamp 1681620392
transform 1 0 1640 0 1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_232
timestamp 1681620392
transform 1 0 1648 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_233
timestamp 1681620392
transform 1 0 1672 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_234
timestamp 1681620392
transform 1 0 1696 0 1 970
box -8 -3 32 105
use NAND3X1  NAND3X1_91
timestamp 1681620392
transform 1 0 1720 0 1 970
box -8 -3 40 105
use FILL  FILL_999
timestamp 1681620392
transform 1 0 1752 0 1 970
box -8 -3 16 105
use FILL  FILL_1000
timestamp 1681620392
transform 1 0 1760 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_225
timestamp 1681620392
transform 1 0 1768 0 1 970
box -8 -3 104 105
use NAND2X1  NAND2X1_235
timestamp 1681620392
transform 1 0 1864 0 1 970
box -8 -3 32 105
use FILL  FILL_1001
timestamp 1681620392
transform 1 0 1888 0 1 970
box -8 -3 16 105
use FILL  FILL_1002
timestamp 1681620392
transform 1 0 1896 0 1 970
box -8 -3 16 105
use FILL  FILL_1009
timestamp 1681620392
transform 1 0 1904 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_226
timestamp 1681620392
transform 1 0 1912 0 1 970
box -8 -3 104 105
use FILL  FILL_1011
timestamp 1681620392
transform 1 0 2008 0 1 970
box -8 -3 16 105
use INVX2  INVX2_271
timestamp 1681620392
transform 1 0 2016 0 1 970
box -9 -3 26 105
use OAI22X1  OAI22X1_75
timestamp 1681620392
transform 1 0 2032 0 1 970
box -8 -3 46 105
use FILL  FILL_1013
timestamp 1681620392
transform 1 0 2072 0 1 970
box -8 -3 16 105
use FILL  FILL_1014
timestamp 1681620392
transform 1 0 2080 0 1 970
box -8 -3 16 105
use FILL  FILL_1015
timestamp 1681620392
transform 1 0 2088 0 1 970
box -8 -3 16 105
use FILL  FILL_1016
timestamp 1681620392
transform 1 0 2096 0 1 970
box -8 -3 16 105
use INVX2  INVX2_272
timestamp 1681620392
transform 1 0 2104 0 1 970
box -9 -3 26 105
use INVX2  INVX2_273
timestamp 1681620392
transform 1 0 2120 0 1 970
box -9 -3 26 105
use FILL  FILL_1017
timestamp 1681620392
transform 1 0 2136 0 1 970
box -8 -3 16 105
use FILL  FILL_1018
timestamp 1681620392
transform 1 0 2144 0 1 970
box -8 -3 16 105
use FILL  FILL_1019
timestamp 1681620392
transform 1 0 2152 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_235
timestamp 1681620392
transform 1 0 2160 0 1 970
box -8 -3 34 105
use FILL  FILL_1020
timestamp 1681620392
transform 1 0 2192 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_228
timestamp 1681620392
transform 1 0 2200 0 1 970
box -8 -3 104 105
use NAND2X1  NAND2X1_238
timestamp 1681620392
transform -1 0 2320 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_239
timestamp 1681620392
transform 1 0 2320 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_240
timestamp 1681620392
transform 1 0 2344 0 1 970
box -8 -3 32 105
use FILL  FILL_1023
timestamp 1681620392
transform 1 0 2368 0 1 970
box -8 -3 16 105
use FILL  FILL_1025
timestamp 1681620392
transform 1 0 2376 0 1 970
box -8 -3 16 105
use FILL  FILL_1027
timestamp 1681620392
transform 1 0 2384 0 1 970
box -8 -3 16 105
use FILL  FILL_1028
timestamp 1681620392
transform 1 0 2392 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_237
timestamp 1681620392
transform -1 0 2432 0 1 970
box -8 -3 34 105
use FILL  FILL_1029
timestamp 1681620392
transform 1 0 2432 0 1 970
box -8 -3 16 105
use FILL  FILL_1030
timestamp 1681620392
transform 1 0 2440 0 1 970
box -8 -3 16 105
use FILL  FILL_1033
timestamp 1681620392
transform 1 0 2448 0 1 970
box -8 -3 16 105
use FILL  FILL_1035
timestamp 1681620392
transform 1 0 2456 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_231
timestamp 1681620392
transform 1 0 2464 0 1 970
box -8 -3 104 105
use FILL  FILL_1037
timestamp 1681620392
transform 1 0 2560 0 1 970
box -8 -3 16 105
use INVX2  INVX2_275
timestamp 1681620392
transform 1 0 2568 0 1 970
box -9 -3 26 105
use FILL  FILL_1038
timestamp 1681620392
transform 1 0 2584 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_3407
timestamp 1681620392
transform 1 0 2620 0 1 975
box -3 -3 3 3
use OAI22X1  OAI22X1_77
timestamp 1681620392
transform -1 0 2632 0 1 970
box -8 -3 46 105
use FILL  FILL_1039
timestamp 1681620392
transform 1 0 2632 0 1 970
box -8 -3 16 105
use FILL  FILL_1040
timestamp 1681620392
transform 1 0 2640 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_239
timestamp 1681620392
transform 1 0 2648 0 1 970
box -8 -3 34 105
use M3_M2  M3_M2_3408
timestamp 1681620392
transform 1 0 2700 0 1 975
box -3 -3 3 3
use INVX2  INVX2_276
timestamp 1681620392
transform 1 0 2680 0 1 970
box -9 -3 26 105
use FILL  FILL_1041
timestamp 1681620392
transform 1 0 2696 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_241
timestamp 1681620392
transform 1 0 2704 0 1 970
box -8 -3 34 105
use M3_M2  M3_M2_3409
timestamp 1681620392
transform 1 0 2764 0 1 975
box -3 -3 3 3
use OAI21X1  OAI21X1_242
timestamp 1681620392
transform 1 0 2736 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_243
timestamp 1681620392
transform 1 0 2768 0 1 970
box -8 -3 34 105
use INVX2  INVX2_278
timestamp 1681620392
transform -1 0 2816 0 1 970
box -9 -3 26 105
use FILL  FILL_1049
timestamp 1681620392
transform 1 0 2816 0 1 970
box -8 -3 16 105
use FILL  FILL_1050
timestamp 1681620392
transform 1 0 2824 0 1 970
box -8 -3 16 105
use FILL  FILL_1051
timestamp 1681620392
transform 1 0 2832 0 1 970
box -8 -3 16 105
use FILL  FILL_1052
timestamp 1681620392
transform 1 0 2840 0 1 970
box -8 -3 16 105
use FILL  FILL_1054
timestamp 1681620392
transform 1 0 2848 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_244
timestamp 1681620392
transform 1 0 2856 0 1 970
box -8 -3 34 105
use FILL  FILL_1055
timestamp 1681620392
transform 1 0 2888 0 1 970
box -8 -3 16 105
use FILL  FILL_1056
timestamp 1681620392
transform 1 0 2896 0 1 970
box -8 -3 16 105
use FILL  FILL_1057
timestamp 1681620392
transform 1 0 2904 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_3410
timestamp 1681620392
transform 1 0 2924 0 1 975
box -3 -3 3 3
use OAI21X1  OAI21X1_245
timestamp 1681620392
transform 1 0 2912 0 1 970
box -8 -3 34 105
use FILL  FILL_1059
timestamp 1681620392
transform 1 0 2944 0 1 970
box -8 -3 16 105
use FILL  FILL_1060
timestamp 1681620392
transform 1 0 2952 0 1 970
box -8 -3 16 105
use FILL  FILL_1061
timestamp 1681620392
transform 1 0 2960 0 1 970
box -8 -3 16 105
use FILL  FILL_1063
timestamp 1681620392
transform 1 0 2968 0 1 970
box -8 -3 16 105
use FILL  FILL_1064
timestamp 1681620392
transform 1 0 2976 0 1 970
box -8 -3 16 105
use INVX2  INVX2_280
timestamp 1681620392
transform 1 0 2984 0 1 970
box -9 -3 26 105
use FILL  FILL_1065
timestamp 1681620392
transform 1 0 3000 0 1 970
box -8 -3 16 105
use FILL  FILL_1068
timestamp 1681620392
transform 1 0 3008 0 1 970
box -8 -3 16 105
use Project_Top_VIA0  Project_Top_VIA0_41
timestamp 1681620392
transform 1 0 3043 0 1 970
box -10 -3 10 3
use M3_M2  M3_M2_3446
timestamp 1681620392
transform 1 0 132 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3447
timestamp 1681620392
transform 1 0 188 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_3939
timestamp 1681620392
transform 1 0 84 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3940
timestamp 1681620392
transform 1 0 172 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3941
timestamp 1681620392
transform 1 0 188 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3492
timestamp 1681620392
transform 1 0 84 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4025
timestamp 1681620392
transform 1 0 132 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4026
timestamp 1681620392
transform 1 0 164 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4027
timestamp 1681620392
transform 1 0 180 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4028
timestamp 1681620392
transform 1 0 196 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3519
timestamp 1681620392
transform 1 0 180 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_3936
timestamp 1681620392
transform 1 0 220 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_3942
timestamp 1681620392
transform 1 0 212 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3520
timestamp 1681620392
transform 1 0 228 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3493
timestamp 1681620392
transform 1 0 244 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4029
timestamp 1681620392
transform 1 0 252 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3943
timestamp 1681620392
transform 1 0 276 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3944
timestamp 1681620392
transform 1 0 284 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3494
timestamp 1681620392
transform 1 0 316 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4030
timestamp 1681620392
transform 1 0 324 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4113
timestamp 1681620392
transform 1 0 316 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3945
timestamp 1681620392
transform 1 0 348 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4031
timestamp 1681620392
transform 1 0 340 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3495
timestamp 1681620392
transform 1 0 348 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3544
timestamp 1681620392
transform 1 0 332 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3562
timestamp 1681620392
transform 1 0 324 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3473
timestamp 1681620392
transform 1 0 364 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_3946
timestamp 1681620392
transform 1 0 372 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4032
timestamp 1681620392
transform 1 0 364 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4033
timestamp 1681620392
transform 1 0 380 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4034
timestamp 1681620392
transform 1 0 388 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4114
timestamp 1681620392
transform 1 0 364 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_3521
timestamp 1681620392
transform 1 0 380 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_4115
timestamp 1681620392
transform 1 0 388 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4116
timestamp 1681620392
transform 1 0 396 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_3545
timestamp 1681620392
transform 1 0 364 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_3947
timestamp 1681620392
transform 1 0 412 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3496
timestamp 1681620392
transform 1 0 412 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4035
timestamp 1681620392
transform 1 0 420 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4036
timestamp 1681620392
transform 1 0 428 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4117
timestamp 1681620392
transform 1 0 436 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4150
timestamp 1681620392
transform 1 0 444 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_3563
timestamp 1681620392
transform 1 0 444 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_4037
timestamp 1681620392
transform 1 0 460 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3522
timestamp 1681620392
transform 1 0 460 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3429
timestamp 1681620392
transform 1 0 564 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_3948
timestamp 1681620392
transform 1 0 524 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3474
timestamp 1681620392
transform 1 0 548 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3475
timestamp 1681620392
transform 1 0 572 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_4038
timestamp 1681620392
transform 1 0 500 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3497
timestamp 1681620392
transform 1 0 516 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4039
timestamp 1681620392
transform 1 0 532 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4040
timestamp 1681620392
transform 1 0 548 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4118
timestamp 1681620392
transform 1 0 484 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4119
timestamp 1681620392
transform 1 0 492 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_3564
timestamp 1681620392
transform 1 0 484 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3523
timestamp 1681620392
transform 1 0 500 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_4120
timestamp 1681620392
transform 1 0 516 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4151
timestamp 1681620392
transform 1 0 508 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_3949
timestamp 1681620392
transform 1 0 604 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3448
timestamp 1681620392
transform 1 0 644 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_3950
timestamp 1681620392
transform 1 0 628 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3951
timestamp 1681620392
transform 1 0 636 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4041
timestamp 1681620392
transform 1 0 580 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4042
timestamp 1681620392
transform 1 0 604 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4121
timestamp 1681620392
transform 1 0 548 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4122
timestamp 1681620392
transform 1 0 564 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4123
timestamp 1681620392
transform 1 0 572 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4152
timestamp 1681620392
transform 1 0 540 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_4153
timestamp 1681620392
transform 1 0 556 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_3498
timestamp 1681620392
transform 1 0 612 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3499
timestamp 1681620392
transform 1 0 628 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4124
timestamp 1681620392
transform 1 0 596 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4154
timestamp 1681620392
transform 1 0 588 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_3577
timestamp 1681620392
transform 1 0 588 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_4125
timestamp 1681620392
transform 1 0 628 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_3476
timestamp 1681620392
transform 1 0 660 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_4043
timestamp 1681620392
transform 1 0 644 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4044
timestamp 1681620392
transform 1 0 660 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3411
timestamp 1681620392
transform 1 0 740 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3430
timestamp 1681620392
transform 1 0 748 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3449
timestamp 1681620392
transform 1 0 700 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3450
timestamp 1681620392
transform 1 0 724 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3412
timestamp 1681620392
transform 1 0 780 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_3952
timestamp 1681620392
transform 1 0 700 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3953
timestamp 1681620392
transform 1 0 708 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3954
timestamp 1681620392
transform 1 0 724 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3955
timestamp 1681620392
transform 1 0 740 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3956
timestamp 1681620392
transform 1 0 748 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3957
timestamp 1681620392
transform 1 0 764 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3958
timestamp 1681620392
transform 1 0 780 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3959
timestamp 1681620392
transform 1 0 796 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4045
timestamp 1681620392
transform 1 0 700 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4046
timestamp 1681620392
transform 1 0 716 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4047
timestamp 1681620392
transform 1 0 732 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4126
timestamp 1681620392
transform 1 0 660 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4127
timestamp 1681620392
transform 1 0 676 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4128
timestamp 1681620392
transform 1 0 684 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4155
timestamp 1681620392
transform 1 0 652 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_3524
timestamp 1681620392
transform 1 0 700 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3546
timestamp 1681620392
transform 1 0 676 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3578
timestamp 1681620392
transform 1 0 660 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3579
timestamp 1681620392
transform 1 0 684 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3547
timestamp 1681620392
transform 1 0 716 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3565
timestamp 1681620392
transform 1 0 708 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3477
timestamp 1681620392
transform 1 0 820 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3431
timestamp 1681620392
transform 1 0 916 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3432
timestamp 1681620392
transform 1 0 948 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_3960
timestamp 1681620392
transform 1 0 884 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4048
timestamp 1681620392
transform 1 0 756 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4049
timestamp 1681620392
transform 1 0 780 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4050
timestamp 1681620392
transform 1 0 820 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3525
timestamp 1681620392
transform 1 0 756 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3500
timestamp 1681620392
transform 1 0 828 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3478
timestamp 1681620392
transform 1 0 892 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_3961
timestamp 1681620392
transform 1 0 908 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3962
timestamp 1681620392
transform 1 0 916 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3479
timestamp 1681620392
transform 1 0 924 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_3963
timestamp 1681620392
transform 1 0 940 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4051
timestamp 1681620392
transform 1 0 876 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4052
timestamp 1681620392
transform 1 0 892 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3501
timestamp 1681620392
transform 1 0 916 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4053
timestamp 1681620392
transform 1 0 924 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3502
timestamp 1681620392
transform 1 0 940 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4129
timestamp 1681620392
transform 1 0 908 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_3413
timestamp 1681620392
transform 1 0 980 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_3964
timestamp 1681620392
transform 1 0 956 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3480
timestamp 1681620392
transform 1 0 964 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3451
timestamp 1681620392
transform 1 0 1060 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_3965
timestamp 1681620392
transform 1 0 980 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3966
timestamp 1681620392
transform 1 0 996 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4130
timestamp 1681620392
transform 1 0 948 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4131
timestamp 1681620392
transform 1 0 956 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_3566
timestamp 1681620392
transform 1 0 940 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3548
timestamp 1681620392
transform 1 0 956 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3481
timestamp 1681620392
transform 1 0 1020 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3414
timestamp 1681620392
transform 1 0 1100 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3433
timestamp 1681620392
transform 1 0 1108 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3452
timestamp 1681620392
transform 1 0 1108 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_3967
timestamp 1681620392
transform 1 0 1100 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4054
timestamp 1681620392
transform 1 0 980 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4055
timestamp 1681620392
transform 1 0 1020 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4056
timestamp 1681620392
transform 1 0 1076 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4057
timestamp 1681620392
transform 1 0 1092 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3526
timestamp 1681620392
transform 1 0 980 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3549
timestamp 1681620392
transform 1 0 980 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3550
timestamp 1681620392
transform 1 0 1028 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3567
timestamp 1681620392
transform 1 0 972 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3527
timestamp 1681620392
transform 1 0 1092 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_4058
timestamp 1681620392
transform 1 0 1108 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3415
timestamp 1681620392
transform 1 0 1148 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3453
timestamp 1681620392
transform 1 0 1140 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_3968
timestamp 1681620392
transform 1 0 1140 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3969
timestamp 1681620392
transform 1 0 1148 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4059
timestamp 1681620392
transform 1 0 1124 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3528
timestamp 1681620392
transform 1 0 1124 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_4132
timestamp 1681620392
transform 1 0 1140 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4060
timestamp 1681620392
transform 1 0 1156 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4061
timestamp 1681620392
transform 1 0 1164 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3529
timestamp 1681620392
transform 1 0 1164 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3568
timestamp 1681620392
transform 1 0 1156 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_3970
timestamp 1681620392
transform 1 0 1172 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3971
timestamp 1681620392
transform 1 0 1228 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4062
timestamp 1681620392
transform 1 0 1212 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3580
timestamp 1681620392
transform 1 0 1212 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3569
timestamp 1681620392
transform 1 0 1244 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_3972
timestamp 1681620392
transform 1 0 1260 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3973
timestamp 1681620392
transform 1 0 1276 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3482
timestamp 1681620392
transform 1 0 1292 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3454
timestamp 1681620392
transform 1 0 1324 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_3974
timestamp 1681620392
transform 1 0 1324 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3975
timestamp 1681620392
transform 1 0 1332 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4063
timestamp 1681620392
transform 1 0 1300 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4064
timestamp 1681620392
transform 1 0 1316 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4133
timestamp 1681620392
transform 1 0 1292 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_3530
timestamp 1681620392
transform 1 0 1316 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3551
timestamp 1681620392
transform 1 0 1300 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3483
timestamp 1681620392
transform 1 0 1356 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3484
timestamp 1681620392
transform 1 0 1372 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_4065
timestamp 1681620392
transform 1 0 1348 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4066
timestamp 1681620392
transform 1 0 1356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4067
timestamp 1681620392
transform 1 0 1364 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3416
timestamp 1681620392
transform 1 0 1388 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3434
timestamp 1681620392
transform 1 0 1420 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_3976
timestamp 1681620392
transform 1 0 1388 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3977
timestamp 1681620392
transform 1 0 1396 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3978
timestamp 1681620392
transform 1 0 1412 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3979
timestamp 1681620392
transform 1 0 1420 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3980
timestamp 1681620392
transform 1 0 1452 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3981
timestamp 1681620392
transform 1 0 1460 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4068
timestamp 1681620392
transform 1 0 1388 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3503
timestamp 1681620392
transform 1 0 1396 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4069
timestamp 1681620392
transform 1 0 1404 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4070
timestamp 1681620392
transform 1 0 1420 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4071
timestamp 1681620392
transform 1 0 1428 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4072
timestamp 1681620392
transform 1 0 1444 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4073
timestamp 1681620392
transform 1 0 1460 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3552
timestamp 1681620392
transform 1 0 1420 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3570
timestamp 1681620392
transform 1 0 1388 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3571
timestamp 1681620392
transform 1 0 1428 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3581
timestamp 1681620392
transform 1 0 1396 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3553
timestamp 1681620392
transform 1 0 1460 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3417
timestamp 1681620392
transform 1 0 1492 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3418
timestamp 1681620392
transform 1 0 1516 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3435
timestamp 1681620392
transform 1 0 1500 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3455
timestamp 1681620392
transform 1 0 1500 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_3982
timestamp 1681620392
transform 1 0 1508 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3983
timestamp 1681620392
transform 1 0 1524 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4074
timestamp 1681620392
transform 1 0 1484 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4075
timestamp 1681620392
transform 1 0 1500 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4076
timestamp 1681620392
transform 1 0 1516 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3572
timestamp 1681620392
transform 1 0 1476 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3531
timestamp 1681620392
transform 1 0 1524 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3573
timestamp 1681620392
transform 1 0 1516 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3456
timestamp 1681620392
transform 1 0 1556 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_3984
timestamp 1681620392
transform 1 0 1556 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4077
timestamp 1681620392
transform 1 0 1564 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4134
timestamp 1681620392
transform 1 0 1556 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_3554
timestamp 1681620392
transform 1 0 1564 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3436
timestamp 1681620392
transform 1 0 1580 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_3985
timestamp 1681620392
transform 1 0 1580 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4135
timestamp 1681620392
transform 1 0 1580 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4078
timestamp 1681620392
transform 1 0 1596 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3986
timestamp 1681620392
transform 1 0 1612 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4079
timestamp 1681620392
transform 1 0 1620 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4136
timestamp 1681620392
transform 1 0 1612 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_3574
timestamp 1681620392
transform 1 0 1620 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_3987
timestamp 1681620392
transform 1 0 1636 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4080
timestamp 1681620392
transform 1 0 1652 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3988
timestamp 1681620392
transform 1 0 1676 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4081
timestamp 1681620392
transform 1 0 1676 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4137
timestamp 1681620392
transform 1 0 1668 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_3582
timestamp 1681620392
transform 1 0 1668 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_3989
timestamp 1681620392
transform 1 0 1716 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4082
timestamp 1681620392
transform 1 0 1700 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3504
timestamp 1681620392
transform 1 0 1716 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3532
timestamp 1681620392
transform 1 0 1700 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_4138
timestamp 1681620392
transform 1 0 1716 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_3583
timestamp 1681620392
transform 1 0 1684 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3584
timestamp 1681620392
transform 1 0 1716 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_3990
timestamp 1681620392
transform 1 0 1732 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4083
timestamp 1681620392
transform 1 0 1724 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3533
timestamp 1681620392
transform 1 0 1748 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3457
timestamp 1681620392
transform 1 0 1764 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_3991
timestamp 1681620392
transform 1 0 1772 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3485
timestamp 1681620392
transform 1 0 1780 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3458
timestamp 1681620392
transform 1 0 1820 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_3992
timestamp 1681620392
transform 1 0 1788 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3993
timestamp 1681620392
transform 1 0 1796 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3994
timestamp 1681620392
transform 1 0 1812 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3505
timestamp 1681620392
transform 1 0 1764 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4084
timestamp 1681620392
transform 1 0 1780 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3506
timestamp 1681620392
transform 1 0 1788 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4085
timestamp 1681620392
transform 1 0 1804 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4086
timestamp 1681620392
transform 1 0 1820 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4139
timestamp 1681620392
transform 1 0 1756 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_3585
timestamp 1681620392
transform 1 0 1756 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_4140
timestamp 1681620392
transform 1 0 1764 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_3534
timestamp 1681620392
transform 1 0 1780 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3555
timestamp 1681620392
transform 1 0 1772 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3535
timestamp 1681620392
transform 1 0 1804 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3556
timestamp 1681620392
transform 1 0 1796 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3536
timestamp 1681620392
transform 1 0 1844 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_3995
timestamp 1681620392
transform 1 0 1860 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3996
timestamp 1681620392
transform 1 0 1868 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3507
timestamp 1681620392
transform 1 0 1868 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3437
timestamp 1681620392
transform 1 0 1884 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3486
timestamp 1681620392
transform 1 0 1892 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_4087
timestamp 1681620392
transform 1 0 1876 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4088
timestamp 1681620392
transform 1 0 1884 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3537
timestamp 1681620392
transform 1 0 1876 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_4141
timestamp 1681620392
transform 1 0 1892 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_3538
timestamp 1681620392
transform 1 0 1900 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_3997
timestamp 1681620392
transform 1 0 1924 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3487
timestamp 1681620392
transform 1 0 2004 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_4089
timestamp 1681620392
transform 1 0 1948 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4090
timestamp 1681620392
transform 1 0 2004 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3419
timestamp 1681620392
transform 1 0 2020 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3420
timestamp 1681620392
transform 1 0 2060 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3421
timestamp 1681620392
transform 1 0 2084 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3422
timestamp 1681620392
transform 1 0 2124 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3438
timestamp 1681620392
transform 1 0 2116 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3439
timestamp 1681620392
transform 1 0 2132 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3440
timestamp 1681620392
transform 1 0 2148 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3459
timestamp 1681620392
transform 1 0 2076 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3460
timestamp 1681620392
transform 1 0 2132 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_3998
timestamp 1681620392
transform 1 0 2028 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3999
timestamp 1681620392
transform 1 0 2116 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4000
timestamp 1681620392
transform 1 0 2132 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4001
timestamp 1681620392
transform 1 0 2148 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4002
timestamp 1681620392
transform 1 0 2156 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3508
timestamp 1681620392
transform 1 0 2052 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4091
timestamp 1681620392
transform 1 0 2076 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4092
timestamp 1681620392
transform 1 0 2108 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4093
timestamp 1681620392
transform 1 0 2124 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3557
timestamp 1681620392
transform 1 0 2052 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3575
timestamp 1681620392
transform 1 0 2068 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3509
timestamp 1681620392
transform 1 0 2132 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4094
timestamp 1681620392
transform 1 0 2140 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3558
timestamp 1681620392
transform 1 0 2156 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3576
timestamp 1681620392
transform 1 0 2156 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3461
timestamp 1681620392
transform 1 0 2188 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3462
timestamp 1681620392
transform 1 0 2244 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_4003
timestamp 1681620392
transform 1 0 2188 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4004
timestamp 1681620392
transform 1 0 2204 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4005
timestamp 1681620392
transform 1 0 2220 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3510
timestamp 1681620392
transform 1 0 2204 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4095
timestamp 1681620392
transform 1 0 2244 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3511
timestamp 1681620392
transform 1 0 2292 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4006
timestamp 1681620392
transform 1 0 2324 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4096
timestamp 1681620392
transform 1 0 2300 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4097
timestamp 1681620392
transform 1 0 2316 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4142
timestamp 1681620392
transform 1 0 2188 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4143
timestamp 1681620392
transform 1 0 2308 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_3586
timestamp 1681620392
transform 1 0 2228 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3587
timestamp 1681620392
transform 1 0 2316 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3512
timestamp 1681620392
transform 1 0 2340 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4144
timestamp 1681620392
transform 1 0 2364 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4007
timestamp 1681620392
transform 1 0 2388 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4145
timestamp 1681620392
transform 1 0 2380 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4098
timestamp 1681620392
transform 1 0 2396 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4099
timestamp 1681620392
transform 1 0 2412 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3539
timestamp 1681620392
transform 1 0 2396 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3513
timestamp 1681620392
transform 1 0 2420 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3540
timestamp 1681620392
transform 1 0 2436 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_4146
timestamp 1681620392
transform 1 0 2444 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_3463
timestamp 1681620392
transform 1 0 2476 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_4008
timestamp 1681620392
transform 1 0 2476 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4100
timestamp 1681620392
transform 1 0 2468 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3541
timestamp 1681620392
transform 1 0 2468 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3441
timestamp 1681620392
transform 1 0 2500 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_4009
timestamp 1681620392
transform 1 0 2484 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3488
timestamp 1681620392
transform 1 0 2492 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3442
timestamp 1681620392
transform 1 0 2524 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3443
timestamp 1681620392
transform 1 0 2612 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3464
timestamp 1681620392
transform 1 0 2524 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_4010
timestamp 1681620392
transform 1 0 2508 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4011
timestamp 1681620392
transform 1 0 2524 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3489
timestamp 1681620392
transform 1 0 2548 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3490
timestamp 1681620392
transform 1 0 2604 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_4012
timestamp 1681620392
transform 1 0 2612 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3514
timestamp 1681620392
transform 1 0 2492 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4101
timestamp 1681620392
transform 1 0 2500 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3515
timestamp 1681620392
transform 1 0 2508 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4102
timestamp 1681620392
transform 1 0 2548 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3516
timestamp 1681620392
transform 1 0 2612 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3423
timestamp 1681620392
transform 1 0 2628 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_4013
timestamp 1681620392
transform 1 0 2628 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4103
timestamp 1681620392
transform 1 0 2620 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3424
timestamp 1681620392
transform 1 0 2676 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3465
timestamp 1681620392
transform 1 0 2668 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_4014
timestamp 1681620392
transform 1 0 2652 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4015
timestamp 1681620392
transform 1 0 2668 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4016
timestamp 1681620392
transform 1 0 2676 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4104
timestamp 1681620392
transform 1 0 2660 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3425
timestamp 1681620392
transform 1 0 2708 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3426
timestamp 1681620392
transform 1 0 2740 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3427
timestamp 1681620392
transform 1 0 2804 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3466
timestamp 1681620392
transform 1 0 2740 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3467
timestamp 1681620392
transform 1 0 2756 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3491
timestamp 1681620392
transform 1 0 2716 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_4017
timestamp 1681620392
transform 1 0 2724 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4018
timestamp 1681620392
transform 1 0 2740 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4019
timestamp 1681620392
transform 1 0 2756 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4105
timestamp 1681620392
transform 1 0 2716 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3517
timestamp 1681620392
transform 1 0 2724 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4106
timestamp 1681620392
transform 1 0 2732 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3542
timestamp 1681620392
transform 1 0 2716 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3444
timestamp 1681620392
transform 1 0 2852 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3468
timestamp 1681620392
transform 1 0 2844 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_4107
timestamp 1681620392
transform 1 0 2780 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4108
timestamp 1681620392
transform 1 0 2836 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4020
timestamp 1681620392
transform 1 0 2852 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3428
timestamp 1681620392
transform 1 0 2876 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_4109
timestamp 1681620392
transform 1 0 2876 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4147
timestamp 1681620392
transform 1 0 2868 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_3469
timestamp 1681620392
transform 1 0 2900 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3470
timestamp 1681620392
transform 1 0 2932 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_4021
timestamp 1681620392
transform 1 0 2916 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_3518
timestamp 1681620392
transform 1 0 2892 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_4110
timestamp 1681620392
transform 1 0 2900 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4148
timestamp 1681620392
transform 1 0 2884 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4149
timestamp 1681620392
transform 1 0 2900 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_3559
timestamp 1681620392
transform 1 0 2876 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_4156
timestamp 1681620392
transform 1 0 2892 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_3560
timestamp 1681620392
transform 1 0 2900 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3445
timestamp 1681620392
transform 1 0 2956 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_4022
timestamp 1681620392
transform 1 0 2940 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4023
timestamp 1681620392
transform 1 0 2948 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4111
timestamp 1681620392
transform 1 0 2924 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3471
timestamp 1681620392
transform 1 0 2964 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_4112
timestamp 1681620392
transform 1 0 2964 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_3543
timestamp 1681620392
transform 1 0 2964 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3561
timestamp 1681620392
transform 1 0 2972 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3472
timestamp 1681620392
transform 1 0 2988 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_3937
timestamp 1681620392
transform 1 0 2996 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_3938
timestamp 1681620392
transform 1 0 3012 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_4024
timestamp 1681620392
transform 1 0 3004 0 1 935
box -2 -2 2 2
use Project_Top_VIA0  Project_Top_VIA0_42
timestamp 1681620392
transform 1 0 24 0 1 870
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_218
timestamp 1681620392
transform 1 0 72 0 -1 970
box -8 -3 104 105
use OAI22X1  OAI22X1_71
timestamp 1681620392
transform -1 0 208 0 -1 970
box -8 -3 46 105
use FILL  FILL_932
timestamp 1681620392
transform 1 0 208 0 -1 970
box -8 -3 16 105
use FILL  FILL_933
timestamp 1681620392
transform 1 0 216 0 -1 970
box -8 -3 16 105
use FILL  FILL_934
timestamp 1681620392
transform 1 0 224 0 -1 970
box -8 -3 16 105
use NOR2X1  NOR2X1_76
timestamp 1681620392
transform 1 0 232 0 -1 970
box -8 -3 32 105
use FILL  FILL_939
timestamp 1681620392
transform 1 0 256 0 -1 970
box -8 -3 16 105
use FILL  FILL_940
timestamp 1681620392
transform 1 0 264 0 -1 970
box -8 -3 16 105
use FILL  FILL_941
timestamp 1681620392
transform 1 0 272 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_219
timestamp 1681620392
transform 1 0 280 0 -1 970
box -8 -3 32 105
use FILL  FILL_942
timestamp 1681620392
transform 1 0 304 0 -1 970
box -8 -3 16 105
use FILL  FILL_943
timestamp 1681620392
transform 1 0 312 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_254
timestamp 1681620392
transform 1 0 320 0 -1 970
box -9 -3 26 105
use FILL  FILL_944
timestamp 1681620392
transform 1 0 336 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_223
timestamp 1681620392
transform 1 0 344 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_224
timestamp 1681620392
transform 1 0 368 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_225
timestamp 1681620392
transform -1 0 416 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_226
timestamp 1681620392
transform 1 0 416 0 -1 970
box -8 -3 32 105
use FILL  FILL_945
timestamp 1681620392
transform 1 0 440 0 -1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_85
timestamp 1681620392
transform 1 0 448 0 -1 970
box -8 -3 40 105
use FILL  FILL_963
timestamp 1681620392
transform 1 0 480 0 -1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_87
timestamp 1681620392
transform 1 0 488 0 -1 970
box -8 -3 40 105
use INVX2  INVX2_261
timestamp 1681620392
transform 1 0 520 0 -1 970
box -9 -3 26 105
use NAND3X1  NAND3X1_88
timestamp 1681620392
transform 1 0 536 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_89
timestamp 1681620392
transform 1 0 568 0 -1 970
box -8 -3 40 105
use M3_M2  M3_M2_3588
timestamp 1681620392
transform 1 0 628 0 1 875
box -3 -3 3 3
use OAI21X1  OAI21X1_225
timestamp 1681620392
transform 1 0 600 0 -1 970
box -8 -3 34 105
use INVX2  INVX2_262
timestamp 1681620392
transform 1 0 632 0 -1 970
box -9 -3 26 105
use NAND3X1  NAND3X1_90
timestamp 1681620392
transform 1 0 648 0 -1 970
box -8 -3 40 105
use NAND2X1  NAND2X1_227
timestamp 1681620392
transform -1 0 704 0 -1 970
box -8 -3 32 105
use M3_M2  M3_M2_3589
timestamp 1681620392
transform 1 0 724 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_3590
timestamp 1681620392
transform 1 0 740 0 1 875
box -3 -3 3 3
use OAI22X1  OAI22X1_72
timestamp 1681620392
transform -1 0 744 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_73
timestamp 1681620392
transform -1 0 784 0 -1 970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_222
timestamp 1681620392
transform 1 0 784 0 -1 970
box -8 -3 104 105
use OAI21X1  OAI21X1_226
timestamp 1681620392
transform 1 0 880 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_227
timestamp 1681620392
transform 1 0 912 0 -1 970
box -8 -3 34 105
use FILL  FILL_964
timestamp 1681620392
transform 1 0 944 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_228
timestamp 1681620392
transform -1 0 984 0 -1 970
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_223
timestamp 1681620392
transform 1 0 984 0 -1 970
box -8 -3 104 105
use INVX2  INVX2_263
timestamp 1681620392
transform 1 0 1080 0 -1 970
box -9 -3 26 105
use FILL  FILL_965
timestamp 1681620392
transform 1 0 1096 0 -1 970
box -8 -3 16 105
use FILL  FILL_966
timestamp 1681620392
transform 1 0 1104 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_229
timestamp 1681620392
transform 1 0 1112 0 -1 970
box -8 -3 34 105
use INVX2  INVX2_264
timestamp 1681620392
transform 1 0 1144 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_265
timestamp 1681620392
transform -1 0 1176 0 -1 970
box -9 -3 26 105
use FILL  FILL_967
timestamp 1681620392
transform 1 0 1176 0 -1 970
box -8 -3 16 105
use FILL  FILL_968
timestamp 1681620392
transform 1 0 1184 0 -1 970
box -8 -3 16 105
use FILL  FILL_969
timestamp 1681620392
transform 1 0 1192 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_230
timestamp 1681620392
transform 1 0 1200 0 -1 970
box -8 -3 34 105
use FILL  FILL_970
timestamp 1681620392
transform 1 0 1232 0 -1 970
box -8 -3 16 105
use FILL  FILL_971
timestamp 1681620392
transform 1 0 1240 0 -1 970
box -8 -3 16 105
use FILL  FILL_972
timestamp 1681620392
transform 1 0 1248 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_228
timestamp 1681620392
transform 1 0 1256 0 -1 970
box -8 -3 32 105
use FILL  FILL_973
timestamp 1681620392
transform 1 0 1280 0 -1 970
box -8 -3 16 105
use FILL  FILL_975
timestamp 1681620392
transform 1 0 1288 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_37
timestamp 1681620392
transform 1 0 1296 0 -1 970
box -8 -3 46 105
use FILL  FILL_977
timestamp 1681620392
transform 1 0 1336 0 -1 970
box -8 -3 16 105
use FILL  FILL_981
timestamp 1681620392
transform 1 0 1344 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_267
timestamp 1681620392
transform -1 0 1368 0 -1 970
box -9 -3 26 105
use FILL  FILL_982
timestamp 1681620392
transform 1 0 1368 0 -1 970
box -8 -3 16 105
use FILL  FILL_983
timestamp 1681620392
transform 1 0 1376 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_38
timestamp 1681620392
transform -1 0 1424 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_39
timestamp 1681620392
transform -1 0 1464 0 -1 970
box -8 -3 46 105
use FILL  FILL_984
timestamp 1681620392
transform 1 0 1464 0 -1 970
box -8 -3 16 105
use FILL  FILL_985
timestamp 1681620392
transform 1 0 1472 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_41
timestamp 1681620392
transform 1 0 1480 0 -1 970
box -8 -3 46 105
use FILL  FILL_987
timestamp 1681620392
transform 1 0 1520 0 -1 970
box -8 -3 16 105
use FILL  FILL_989
timestamp 1681620392
transform 1 0 1528 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_229
timestamp 1681620392
transform 1 0 1536 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_230
timestamp 1681620392
transform 1 0 1560 0 -1 970
box -8 -3 32 105
use FILL  FILL_996
timestamp 1681620392
transform 1 0 1584 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_231
timestamp 1681620392
transform 1 0 1592 0 -1 970
box -8 -3 32 105
use INVX2  INVX2_268
timestamp 1681620392
transform 1 0 1616 0 -1 970
box -9 -3 26 105
use FILL  FILL_997
timestamp 1681620392
transform 1 0 1632 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_232
timestamp 1681620392
transform 1 0 1640 0 -1 970
box -8 -3 34 105
use INVX2  INVX2_269
timestamp 1681620392
transform 1 0 1672 0 -1 970
box -9 -3 26 105
use OAI21X1  OAI21X1_233
timestamp 1681620392
transform 1 0 1688 0 -1 970
box -8 -3 34 105
use FILL  FILL_1003
timestamp 1681620392
transform 1 0 1720 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_234
timestamp 1681620392
transform 1 0 1728 0 -1 970
box -8 -3 34 105
use FILL  FILL_1004
timestamp 1681620392
transform 1 0 1760 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_236
timestamp 1681620392
transform -1 0 1792 0 -1 970
box -8 -3 32 105
use OAI22X1  OAI22X1_74
timestamp 1681620392
transform -1 0 1832 0 -1 970
box -8 -3 46 105
use INVX2  INVX2_270
timestamp 1681620392
transform -1 0 1848 0 -1 970
box -9 -3 26 105
use FILL  FILL_1005
timestamp 1681620392
transform 1 0 1848 0 -1 970
box -8 -3 16 105
use FILL  FILL_1006
timestamp 1681620392
transform 1 0 1856 0 -1 970
box -8 -3 16 105
use FILL  FILL_1007
timestamp 1681620392
transform 1 0 1864 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_237
timestamp 1681620392
transform 1 0 1872 0 -1 970
box -8 -3 32 105
use FILL  FILL_1008
timestamp 1681620392
transform 1 0 1896 0 -1 970
box -8 -3 16 105
use FILL  FILL_1010
timestamp 1681620392
transform 1 0 1904 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_227
timestamp 1681620392
transform 1 0 1912 0 -1 970
box -8 -3 104 105
use FILL  FILL_1012
timestamp 1681620392
transform 1 0 2008 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_229
timestamp 1681620392
transform 1 0 2016 0 -1 970
box -8 -3 104 105
use OAI22X1  OAI22X1_76
timestamp 1681620392
transform -1 0 2152 0 -1 970
box -8 -3 46 105
use OAI21X1  OAI21X1_236
timestamp 1681620392
transform 1 0 2152 0 -1 970
box -8 -3 34 105
use NAND2X1  NAND2X1_241
timestamp 1681620392
transform -1 0 2208 0 -1 970
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_230
timestamp 1681620392
transform 1 0 2208 0 -1 970
box -8 -3 104 105
use NAND2X1  NAND2X1_242
timestamp 1681620392
transform -1 0 2328 0 -1 970
box -8 -3 32 105
use FILL  FILL_1021
timestamp 1681620392
transform 1 0 2328 0 -1 970
box -8 -3 16 105
use FILL  FILL_1022
timestamp 1681620392
transform 1 0 2336 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_243
timestamp 1681620392
transform 1 0 2344 0 -1 970
box -8 -3 32 105
use FILL  FILL_1024
timestamp 1681620392
transform 1 0 2368 0 -1 970
box -8 -3 16 105
use FILL  FILL_1026
timestamp 1681620392
transform 1 0 2376 0 -1 970
box -8 -3 16 105
use FILL  FILL_1031
timestamp 1681620392
transform 1 0 2384 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_238
timestamp 1681620392
transform -1 0 2424 0 -1 970
box -8 -3 34 105
use INVX2  INVX2_274
timestamp 1681620392
transform -1 0 2440 0 -1 970
box -9 -3 26 105
use FILL  FILL_1032
timestamp 1681620392
transform 1 0 2440 0 -1 970
box -8 -3 16 105
use FILL  FILL_1034
timestamp 1681620392
transform 1 0 2448 0 -1 970
box -8 -3 16 105
use FILL  FILL_1036
timestamp 1681620392
transform 1 0 2456 0 -1 970
box -8 -3 16 105
use FILL  FILL_1042
timestamp 1681620392
transform 1 0 2464 0 -1 970
box -8 -3 16 105
use FILL  FILL_1043
timestamp 1681620392
transform 1 0 2472 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_240
timestamp 1681620392
transform -1 0 2512 0 -1 970
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_232
timestamp 1681620392
transform 1 0 2512 0 -1 970
box -8 -3 104 105
use INVX2  INVX2_277
timestamp 1681620392
transform 1 0 2608 0 -1 970
box -9 -3 26 105
use FILL  FILL_1044
timestamp 1681620392
transform 1 0 2624 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_78
timestamp 1681620392
transform 1 0 2632 0 -1 970
box -8 -3 46 105
use FILL  FILL_1045
timestamp 1681620392
transform 1 0 2672 0 -1 970
box -8 -3 16 105
use FILL  FILL_1046
timestamp 1681620392
transform 1 0 2680 0 -1 970
box -8 -3 16 105
use FILL  FILL_1047
timestamp 1681620392
transform 1 0 2688 0 -1 970
box -8 -3 16 105
use FILL  FILL_1048
timestamp 1681620392
transform 1 0 2696 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_79
timestamp 1681620392
transform 1 0 2704 0 -1 970
box -8 -3 46 105
use M3_M2  M3_M2_3591
timestamp 1681620392
transform 1 0 2764 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_3592
timestamp 1681620392
transform 1 0 2828 0 1 875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_233
timestamp 1681620392
transform 1 0 2744 0 -1 970
box -8 -3 104 105
use FILL  FILL_1053
timestamp 1681620392
transform 1 0 2840 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_244
timestamp 1681620392
transform 1 0 2848 0 -1 970
box -8 -3 32 105
use FILL  FILL_1058
timestamp 1681620392
transform 1 0 2872 0 -1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_92
timestamp 1681620392
transform -1 0 2912 0 -1 970
box -8 -3 40 105
use OAI21X1  OAI21X1_246
timestamp 1681620392
transform 1 0 2912 0 -1 970
box -8 -3 34 105
use INVX2  INVX2_279
timestamp 1681620392
transform 1 0 2944 0 -1 970
box -9 -3 26 105
use FILL  FILL_1062
timestamp 1681620392
transform 1 0 2960 0 -1 970
box -8 -3 16 105
use FILL  FILL_1066
timestamp 1681620392
transform 1 0 2968 0 -1 970
box -8 -3 16 105
use NOR2X1  NOR2X1_79
timestamp 1681620392
transform -1 0 3000 0 -1 970
box -8 -3 32 105
use FILL  FILL_1067
timestamp 1681620392
transform 1 0 3000 0 -1 970
box -8 -3 16 105
use FILL  FILL_1069
timestamp 1681620392
transform 1 0 3008 0 -1 970
box -8 -3 16 105
use Project_Top_VIA0  Project_Top_VIA0_43
timestamp 1681620392
transform 1 0 3067 0 1 870
box -10 -3 10 3
use M3_M2  M3_M2_3637
timestamp 1681620392
transform 1 0 140 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_4189
timestamp 1681620392
transform 1 0 140 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4190
timestamp 1681620392
transform 1 0 156 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3638
timestamp 1681620392
transform 1 0 196 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_4191
timestamp 1681620392
transform 1 0 180 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3659
timestamp 1681620392
transform 1 0 188 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4192
timestamp 1681620392
transform 1 0 196 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4270
timestamp 1681620392
transform 1 0 132 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4271
timestamp 1681620392
transform 1 0 148 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4272
timestamp 1681620392
transform 1 0 172 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4273
timestamp 1681620392
transform 1 0 188 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3739
timestamp 1681620392
transform 1 0 132 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3690
timestamp 1681620392
transform 1 0 196 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_4193
timestamp 1681620392
transform 1 0 244 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4194
timestamp 1681620392
transform 1 0 300 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4274
timestamp 1681620392
transform 1 0 204 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4275
timestamp 1681620392
transform 1 0 220 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3710
timestamp 1681620392
transform 1 0 188 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3711
timestamp 1681620392
transform 1 0 244 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_4344
timestamp 1681620392
transform 1 0 308 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_3740
timestamp 1681620392
transform 1 0 180 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3741
timestamp 1681620392
transform 1 0 204 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_4159
timestamp 1681620392
transform 1 0 332 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4195
timestamp 1681620392
transform 1 0 324 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3660
timestamp 1681620392
transform 1 0 332 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4276
timestamp 1681620392
transform 1 0 332 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3742
timestamp 1681620392
transform 1 0 316 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3619
timestamp 1681620392
transform 1 0 364 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_4196
timestamp 1681620392
transform 1 0 356 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4277
timestamp 1681620392
transform 1 0 348 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4278
timestamp 1681620392
transform 1 0 364 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3743
timestamp 1681620392
transform 1 0 356 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3620
timestamp 1681620392
transform 1 0 412 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_4160
timestamp 1681620392
transform 1 0 388 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_3639
timestamp 1681620392
transform 1 0 396 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_4161
timestamp 1681620392
transform 1 0 404 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4162
timestamp 1681620392
transform 1 0 412 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4197
timestamp 1681620392
transform 1 0 380 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3661
timestamp 1681620392
transform 1 0 388 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4198
timestamp 1681620392
transform 1 0 396 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4279
timestamp 1681620392
transform 1 0 388 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3712
timestamp 1681620392
transform 1 0 380 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3662
timestamp 1681620392
transform 1 0 420 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3744
timestamp 1681620392
transform 1 0 404 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3621
timestamp 1681620392
transform 1 0 436 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_4199
timestamp 1681620392
transform 1 0 436 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4200
timestamp 1681620392
transform 1 0 444 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4280
timestamp 1681620392
transform 1 0 436 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3713
timestamp 1681620392
transform 1 0 428 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3603
timestamp 1681620392
transform 1 0 476 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3622
timestamp 1681620392
transform 1 0 476 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_4201
timestamp 1681620392
transform 1 0 468 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3691
timestamp 1681620392
transform 1 0 468 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_4281
timestamp 1681620392
transform 1 0 476 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4345
timestamp 1681620392
transform 1 0 468 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_3640
timestamp 1681620392
transform 1 0 500 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_4163
timestamp 1681620392
transform 1 0 524 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4202
timestamp 1681620392
transform 1 0 500 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4203
timestamp 1681620392
transform 1 0 516 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3663
timestamp 1681620392
transform 1 0 524 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3692
timestamp 1681620392
transform 1 0 516 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3745
timestamp 1681620392
transform 1 0 516 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_4164
timestamp 1681620392
transform 1 0 548 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_3641
timestamp 1681620392
transform 1 0 564 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_4204
timestamp 1681620392
transform 1 0 564 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3664
timestamp 1681620392
transform 1 0 572 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4205
timestamp 1681620392
transform 1 0 580 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3665
timestamp 1681620392
transform 1 0 588 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4282
timestamp 1681620392
transform 1 0 564 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4283
timestamp 1681620392
transform 1 0 572 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3693
timestamp 1681620392
transform 1 0 588 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3714
timestamp 1681620392
transform 1 0 564 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3623
timestamp 1681620392
transform 1 0 604 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3604
timestamp 1681620392
transform 1 0 620 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_4157
timestamp 1681620392
transform 1 0 628 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_4165
timestamp 1681620392
transform 1 0 612 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4206
timestamp 1681620392
transform 1 0 604 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3746
timestamp 1681620392
transform 1 0 596 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3666
timestamp 1681620392
transform 1 0 612 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3624
timestamp 1681620392
transform 1 0 684 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_4166
timestamp 1681620392
transform 1 0 636 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4207
timestamp 1681620392
transform 1 0 620 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3642
timestamp 1681620392
transform 1 0 668 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_4167
timestamp 1681620392
transform 1 0 684 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4284
timestamp 1681620392
transform 1 0 644 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3715
timestamp 1681620392
transform 1 0 628 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3747
timestamp 1681620392
transform 1 0 644 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_4208
timestamp 1681620392
transform 1 0 668 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3605
timestamp 1681620392
transform 1 0 708 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3667
timestamp 1681620392
transform 1 0 700 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4209
timestamp 1681620392
transform 1 0 708 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4285
timestamp 1681620392
transform 1 0 700 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4286
timestamp 1681620392
transform 1 0 708 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4168
timestamp 1681620392
transform 1 0 732 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_3643
timestamp 1681620392
transform 1 0 780 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3644
timestamp 1681620392
transform 1 0 836 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3668
timestamp 1681620392
transform 1 0 732 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4210
timestamp 1681620392
transform 1 0 772 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3669
timestamp 1681620392
transform 1 0 796 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4211
timestamp 1681620392
transform 1 0 828 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4212
timestamp 1681620392
transform 1 0 836 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4287
timestamp 1681620392
transform 1 0 732 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4288
timestamp 1681620392
transform 1 0 748 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3748
timestamp 1681620392
transform 1 0 732 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_4169
timestamp 1681620392
transform 1 0 852 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4289
timestamp 1681620392
transform 1 0 844 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3694
timestamp 1681620392
transform 1 0 852 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_4290
timestamp 1681620392
transform 1 0 876 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3716
timestamp 1681620392
transform 1 0 876 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_4213
timestamp 1681620392
transform 1 0 924 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4214
timestamp 1681620392
transform 1 0 956 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4291
timestamp 1681620392
transform 1 0 900 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3670
timestamp 1681620392
transform 1 0 1004 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4292
timestamp 1681620392
transform 1 0 1004 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3717
timestamp 1681620392
transform 1 0 956 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3645
timestamp 1681620392
transform 1 0 1028 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_4215
timestamp 1681620392
transform 1 0 1028 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4346
timestamp 1681620392
transform 1 0 1020 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_3749
timestamp 1681620392
transform 1 0 1020 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_4216
timestamp 1681620392
transform 1 0 1052 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3625
timestamp 1681620392
transform 1 0 1084 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3626
timestamp 1681620392
transform 1 0 1132 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3646
timestamp 1681620392
transform 1 0 1116 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_4217
timestamp 1681620392
transform 1 0 1084 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4218
timestamp 1681620392
transform 1 0 1116 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3671
timestamp 1681620392
transform 1 0 1164 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4293
timestamp 1681620392
transform 1 0 1164 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3750
timestamp 1681620392
transform 1 0 1164 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_4294
timestamp 1681620392
transform 1 0 1180 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4170
timestamp 1681620392
transform 1 0 1212 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_3672
timestamp 1681620392
transform 1 0 1212 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4171
timestamp 1681620392
transform 1 0 1244 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4219
timestamp 1681620392
transform 1 0 1244 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4295
timestamp 1681620392
transform 1 0 1220 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3695
timestamp 1681620392
transform 1 0 1236 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3673
timestamp 1681620392
transform 1 0 1292 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4220
timestamp 1681620392
transform 1 0 1300 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4296
timestamp 1681620392
transform 1 0 1244 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4297
timestamp 1681620392
transform 1 0 1252 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4298
timestamp 1681620392
transform 1 0 1276 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3718
timestamp 1681620392
transform 1 0 1244 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_4347
timestamp 1681620392
transform 1 0 1284 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_3751
timestamp 1681620392
transform 1 0 1276 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_4299
timestamp 1681620392
transform 1 0 1308 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4172
timestamp 1681620392
transform 1 0 1372 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4221
timestamp 1681620392
transform 1 0 1348 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4348
timestamp 1681620392
transform 1 0 1340 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_3719
timestamp 1681620392
transform 1 0 1348 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3647
timestamp 1681620392
transform 1 0 1396 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3674
timestamp 1681620392
transform 1 0 1388 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3612
timestamp 1681620392
transform 1 0 1420 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_4173
timestamp 1681620392
transform 1 0 1428 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4174
timestamp 1681620392
transform 1 0 1436 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4222
timestamp 1681620392
transform 1 0 1396 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4223
timestamp 1681620392
transform 1 0 1412 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4224
timestamp 1681620392
transform 1 0 1420 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4300
timestamp 1681620392
transform 1 0 1380 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4301
timestamp 1681620392
transform 1 0 1404 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4175
timestamp 1681620392
transform 1 0 1460 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_3648
timestamp 1681620392
transform 1 0 1484 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_4225
timestamp 1681620392
transform 1 0 1460 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3675
timestamp 1681620392
transform 1 0 1468 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3593
timestamp 1681620392
transform 1 0 1676 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3627
timestamp 1681620392
transform 1 0 1540 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3628
timestamp 1681620392
transform 1 0 1612 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_4226
timestamp 1681620392
transform 1 0 1476 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4227
timestamp 1681620392
transform 1 0 1484 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4228
timestamp 1681620392
transform 1 0 1508 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4229
timestamp 1681620392
transform 1 0 1524 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4230
timestamp 1681620392
transform 1 0 1556 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4302
timestamp 1681620392
transform 1 0 1452 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3696
timestamp 1681620392
transform 1 0 1460 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3697
timestamp 1681620392
transform 1 0 1476 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_4303
timestamp 1681620392
transform 1 0 1484 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4304
timestamp 1681620392
transform 1 0 1500 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4305
timestamp 1681620392
transform 1 0 1516 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4306
timestamp 1681620392
transform 1 0 1604 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3720
timestamp 1681620392
transform 1 0 1500 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3721
timestamp 1681620392
transform 1 0 1556 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3722
timestamp 1681620392
transform 1 0 1604 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_4231
timestamp 1681620392
transform 1 0 1660 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4307
timestamp 1681620392
transform 1 0 1628 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3723
timestamp 1681620392
transform 1 0 1628 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3724
timestamp 1681620392
transform 1 0 1660 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3594
timestamp 1681620392
transform 1 0 1724 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3613
timestamp 1681620392
transform 1 0 1748 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3649
timestamp 1681620392
transform 1 0 1724 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3650
timestamp 1681620392
transform 1 0 1756 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_4176
timestamp 1681620392
transform 1 0 1764 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4232
timestamp 1681620392
transform 1 0 1716 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4233
timestamp 1681620392
transform 1 0 1724 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4234
timestamp 1681620392
transform 1 0 1732 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4235
timestamp 1681620392
transform 1 0 1748 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4308
timestamp 1681620392
transform 1 0 1740 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4309
timestamp 1681620392
transform 1 0 1756 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3725
timestamp 1681620392
transform 1 0 1740 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3752
timestamp 1681620392
transform 1 0 1748 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_4236
timestamp 1681620392
transform 1 0 1780 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4237
timestamp 1681620392
transform 1 0 1796 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4238
timestamp 1681620392
transform 1 0 1804 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4239
timestamp 1681620392
transform 1 0 1860 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4310
timestamp 1681620392
transform 1 0 1788 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3676
timestamp 1681620392
transform 1 0 1884 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4240
timestamp 1681620392
transform 1 0 1900 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4311
timestamp 1681620392
transform 1 0 1884 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4312
timestamp 1681620392
transform 1 0 1900 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3726
timestamp 1681620392
transform 1 0 1812 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3727
timestamp 1681620392
transform 1 0 1868 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3753
timestamp 1681620392
transform 1 0 1852 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3614
timestamp 1681620392
transform 1 0 1932 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_4177
timestamp 1681620392
transform 1 0 1932 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4313
timestamp 1681620392
transform 1 0 1932 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3615
timestamp 1681620392
transform 1 0 1964 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3629
timestamp 1681620392
transform 1 0 1972 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_4178
timestamp 1681620392
transform 1 0 1980 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4314
timestamp 1681620392
transform 1 0 1972 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3606
timestamp 1681620392
transform 1 0 2076 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3616
timestamp 1681620392
transform 1 0 2044 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3630
timestamp 1681620392
transform 1 0 2004 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3651
timestamp 1681620392
transform 1 0 1996 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_4241
timestamp 1681620392
transform 1 0 1988 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3652
timestamp 1681620392
transform 1 0 2092 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3677
timestamp 1681620392
transform 1 0 2012 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4242
timestamp 1681620392
transform 1 0 2036 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3678
timestamp 1681620392
transform 1 0 2084 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4243
timestamp 1681620392
transform 1 0 2092 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4315
timestamp 1681620392
transform 1 0 1996 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4316
timestamp 1681620392
transform 1 0 2012 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3728
timestamp 1681620392
transform 1 0 1988 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3754
timestamp 1681620392
transform 1 0 1988 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3698
timestamp 1681620392
transform 1 0 2076 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_4317
timestamp 1681620392
transform 1 0 2100 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3729
timestamp 1681620392
transform 1 0 2012 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3730
timestamp 1681620392
transform 1 0 2100 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3755
timestamp 1681620392
transform 1 0 2044 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3607
timestamp 1681620392
transform 1 0 2172 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3617
timestamp 1681620392
transform 1 0 2164 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_4244
timestamp 1681620392
transform 1 0 2116 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3679
timestamp 1681620392
transform 1 0 2124 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4245
timestamp 1681620392
transform 1 0 2132 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3680
timestamp 1681620392
transform 1 0 2148 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4246
timestamp 1681620392
transform 1 0 2156 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3699
timestamp 1681620392
transform 1 0 2116 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_4318
timestamp 1681620392
transform 1 0 2124 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3700
timestamp 1681620392
transform 1 0 2132 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_4319
timestamp 1681620392
transform 1 0 2140 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4320
timestamp 1681620392
transform 1 0 2148 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4321
timestamp 1681620392
transform 1 0 2164 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3701
timestamp 1681620392
transform 1 0 2172 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_4179
timestamp 1681620392
transform 1 0 2228 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_3681
timestamp 1681620392
transform 1 0 2196 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3682
timestamp 1681620392
transform 1 0 2220 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4322
timestamp 1681620392
transform 1 0 2180 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4323
timestamp 1681620392
transform 1 0 2188 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4324
timestamp 1681620392
transform 1 0 2204 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3731
timestamp 1681620392
transform 1 0 2148 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3756
timestamp 1681620392
transform 1 0 2140 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3757
timestamp 1681620392
transform 1 0 2180 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3758
timestamp 1681620392
transform 1 0 2204 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3683
timestamp 1681620392
transform 1 0 2244 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3631
timestamp 1681620392
transform 1 0 2332 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_4247
timestamp 1681620392
transform 1 0 2268 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4248
timestamp 1681620392
transform 1 0 2324 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4325
timestamp 1681620392
transform 1 0 2228 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4326
timestamp 1681620392
transform 1 0 2244 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3732
timestamp 1681620392
transform 1 0 2228 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3733
timestamp 1681620392
transform 1 0 2268 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3759
timestamp 1681620392
transform 1 0 2244 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3760
timestamp 1681620392
transform 1 0 2284 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_4327
timestamp 1681620392
transform 1 0 2332 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3595
timestamp 1681620392
transform 1 0 2348 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3596
timestamp 1681620392
transform 1 0 2380 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3608
timestamp 1681620392
transform 1 0 2364 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3618
timestamp 1681620392
transform 1 0 2372 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3653
timestamp 1681620392
transform 1 0 2356 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3609
timestamp 1681620392
transform 1 0 2436 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3610
timestamp 1681620392
transform 1 0 2460 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3632
timestamp 1681620392
transform 1 0 2388 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3633
timestamp 1681620392
transform 1 0 2428 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_4180
timestamp 1681620392
transform 1 0 2364 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_3702
timestamp 1681620392
transform 1 0 2348 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3654
timestamp 1681620392
transform 1 0 2380 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_4181
timestamp 1681620392
transform 1 0 2388 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4249
timestamp 1681620392
transform 1 0 2372 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4250
timestamp 1681620392
transform 1 0 2380 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3684
timestamp 1681620392
transform 1 0 2388 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4182
timestamp 1681620392
transform 1 0 2492 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4251
timestamp 1681620392
transform 1 0 2428 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4252
timestamp 1681620392
transform 1 0 2484 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4328
timestamp 1681620392
transform 1 0 2364 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3761
timestamp 1681620392
transform 1 0 2356 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3703
timestamp 1681620392
transform 1 0 2380 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3685
timestamp 1681620392
transform 1 0 2492 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4329
timestamp 1681620392
transform 1 0 2404 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4330
timestamp 1681620392
transform 1 0 2492 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3762
timestamp 1681620392
transform 1 0 2396 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3611
timestamp 1681620392
transform 1 0 2516 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3655
timestamp 1681620392
transform 1 0 2524 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_4183
timestamp 1681620392
transform 1 0 2532 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4253
timestamp 1681620392
transform 1 0 2516 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4331
timestamp 1681620392
transform 1 0 2524 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4254
timestamp 1681620392
transform 1 0 2548 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4255
timestamp 1681620392
transform 1 0 2564 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4332
timestamp 1681620392
transform 1 0 2548 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3704
timestamp 1681620392
transform 1 0 2556 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3597
timestamp 1681620392
transform 1 0 2604 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3598
timestamp 1681620392
transform 1 0 2660 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3686
timestamp 1681620392
transform 1 0 2588 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4256
timestamp 1681620392
transform 1 0 2612 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3687
timestamp 1681620392
transform 1 0 2620 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4257
timestamp 1681620392
transform 1 0 2668 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4258
timestamp 1681620392
transform 1 0 2676 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4333
timestamp 1681620392
transform 1 0 2572 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4334
timestamp 1681620392
transform 1 0 2588 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3705
timestamp 1681620392
transform 1 0 2612 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3734
timestamp 1681620392
transform 1 0 2572 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3735
timestamp 1681620392
transform 1 0 2676 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3763
timestamp 1681620392
transform 1 0 2668 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3706
timestamp 1681620392
transform 1 0 2692 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_4259
timestamp 1681620392
transform 1 0 2700 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4335
timestamp 1681620392
transform 1 0 2700 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3764
timestamp 1681620392
transform 1 0 2700 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3634
timestamp 1681620392
transform 1 0 2748 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3656
timestamp 1681620392
transform 1 0 2732 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_4184
timestamp 1681620392
transform 1 0 2748 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4260
timestamp 1681620392
transform 1 0 2732 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4336
timestamp 1681620392
transform 1 0 2724 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3707
timestamp 1681620392
transform 1 0 2740 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_4349
timestamp 1681620392
transform 1 0 2756 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_4261
timestamp 1681620392
transform 1 0 2780 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4350
timestamp 1681620392
transform 1 0 2804 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_4262
timestamp 1681620392
transform 1 0 2820 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4337
timestamp 1681620392
transform 1 0 2836 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4338
timestamp 1681620392
transform 1 0 2844 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3765
timestamp 1681620392
transform 1 0 2844 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_4185
timestamp 1681620392
transform 1 0 2860 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_3599
timestamp 1681620392
transform 1 0 2892 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3600
timestamp 1681620392
transform 1 0 2916 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3635
timestamp 1681620392
transform 1 0 2900 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_4158
timestamp 1681620392
transform 1 0 2916 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_4186
timestamp 1681620392
transform 1 0 2892 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4263
timestamp 1681620392
transform 1 0 2860 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4264
timestamp 1681620392
transform 1 0 2868 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4265
timestamp 1681620392
transform 1 0 2876 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4339
timestamp 1681620392
transform 1 0 2868 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3736
timestamp 1681620392
transform 1 0 2860 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3766
timestamp 1681620392
transform 1 0 2868 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3688
timestamp 1681620392
transform 1 0 2892 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3636
timestamp 1681620392
transform 1 0 2948 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_4187
timestamp 1681620392
transform 1 0 2916 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_3657
timestamp 1681620392
transform 1 0 2924 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3601
timestamp 1681620392
transform 1 0 2964 0 1 865
box -3 -3 3 3
use M2_M1  M2_M1_4188
timestamp 1681620392
transform 1 0 2940 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_3658
timestamp 1681620392
transform 1 0 2956 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_4266
timestamp 1681620392
transform 1 0 2900 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4267
timestamp 1681620392
transform 1 0 2908 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4268
timestamp 1681620392
transform 1 0 2924 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3689
timestamp 1681620392
transform 1 0 2940 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_4340
timestamp 1681620392
transform 1 0 2900 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3708
timestamp 1681620392
transform 1 0 2924 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3709
timestamp 1681620392
transform 1 0 2940 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_4341
timestamp 1681620392
transform 1 0 2948 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4342
timestamp 1681620392
transform 1 0 2956 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_3737
timestamp 1681620392
transform 1 0 2900 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3738
timestamp 1681620392
transform 1 0 2916 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3767
timestamp 1681620392
transform 1 0 2924 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_4343
timestamp 1681620392
transform 1 0 2972 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4351
timestamp 1681620392
transform 1 0 2964 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_4269
timestamp 1681620392
transform 1 0 2980 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_3602
timestamp 1681620392
transform 1 0 2996 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3768
timestamp 1681620392
transform 1 0 2988 0 1 785
box -3 -3 3 3
use Project_Top_VIA0  Project_Top_VIA0_44
timestamp 1681620392
transform 1 0 48 0 1 770
box -10 -3 10 3
use FILL  FILL_1070
timestamp 1681620392
transform 1 0 72 0 1 770
box -8 -3 16 105
use FILL  FILL_1071
timestamp 1681620392
transform 1 0 80 0 1 770
box -8 -3 16 105
use FILL  FILL_1072
timestamp 1681620392
transform 1 0 88 0 1 770
box -8 -3 16 105
use FILL  FILL_1073
timestamp 1681620392
transform 1 0 96 0 1 770
box -8 -3 16 105
use FILL  FILL_1074
timestamp 1681620392
transform 1 0 104 0 1 770
box -8 -3 16 105
use FILL  FILL_1075
timestamp 1681620392
transform 1 0 112 0 1 770
box -8 -3 16 105
use FILL  FILL_1076
timestamp 1681620392
transform 1 0 120 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_80
timestamp 1681620392
transform 1 0 128 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_81
timestamp 1681620392
transform -1 0 208 0 1 770
box -8 -3 46 105
use M3_M2  M3_M2_3769
timestamp 1681620392
transform 1 0 252 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3770
timestamp 1681620392
transform 1 0 308 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_234
timestamp 1681620392
transform 1 0 208 0 1 770
box -8 -3 104 105
use NOR2X1  NOR2X1_80
timestamp 1681620392
transform 1 0 304 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_245
timestamp 1681620392
transform -1 0 352 0 1 770
box -8 -3 32 105
use M3_M2  M3_M2_3771
timestamp 1681620392
transform 1 0 364 0 1 775
box -3 -3 3 3
use FILL  FILL_1077
timestamp 1681620392
transform 1 0 352 0 1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_246
timestamp 1681620392
transform 1 0 360 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_247
timestamp 1681620392
transform 1 0 384 0 1 770
box -8 -3 32 105
use M3_M2  M3_M2_3772
timestamp 1681620392
transform 1 0 436 0 1 775
box -3 -3 3 3
use NAND2X1  NAND2X1_248
timestamp 1681620392
transform -1 0 432 0 1 770
box -8 -3 32 105
use FILL  FILL_1078
timestamp 1681620392
transform 1 0 432 0 1 770
box -8 -3 16 105
use AOI21X1  AOI21X1_26
timestamp 1681620392
transform 1 0 440 0 1 770
box -7 -3 39 105
use FILL  FILL_1079
timestamp 1681620392
transform 1 0 472 0 1 770
box -8 -3 16 105
use FILL  FILL_1085
timestamp 1681620392
transform 1 0 480 0 1 770
box -8 -3 16 105
use AND2X2  AND2X2_23
timestamp 1681620392
transform 1 0 488 0 1 770
box -8 -3 40 105
use FILL  FILL_1087
timestamp 1681620392
transform 1 0 520 0 1 770
box -8 -3 16 105
use FILL  FILL_1088
timestamp 1681620392
transform 1 0 528 0 1 770
box -8 -3 16 105
use FILL  FILL_1089
timestamp 1681620392
transform 1 0 536 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_3773
timestamp 1681620392
transform 1 0 572 0 1 775
box -3 -3 3 3
use NAND2X1  NAND2X1_249
timestamp 1681620392
transform -1 0 568 0 1 770
box -8 -3 32 105
use AND2X2  AND2X2_24
timestamp 1681620392
transform 1 0 568 0 1 770
box -8 -3 40 105
use M3_M2  M3_M2_3774
timestamp 1681620392
transform 1 0 612 0 1 775
box -3 -3 3 3
use FILL  FILL_1090
timestamp 1681620392
transform 1 0 600 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_3775
timestamp 1681620392
transform 1 0 628 0 1 775
box -3 -3 3 3
use NAND3X1  NAND3X1_94
timestamp 1681620392
transform 1 0 608 0 1 770
box -8 -3 40 105
use INVX2  INVX2_285
timestamp 1681620392
transform 1 0 640 0 1 770
box -9 -3 26 105
use OAI21X1  OAI21X1_247
timestamp 1681620392
transform 1 0 656 0 1 770
box -8 -3 34 105
use FILL  FILL_1091
timestamp 1681620392
transform 1 0 688 0 1 770
box -8 -3 16 105
use FILL  FILL_1092
timestamp 1681620392
transform 1 0 696 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_250
timestamp 1681620392
transform 1 0 704 0 1 770
box -8 -3 34 105
use M3_M2  M3_M2_3776
timestamp 1681620392
transform 1 0 748 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3777
timestamp 1681620392
transform 1 0 780 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3778
timestamp 1681620392
transform 1 0 796 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_237
timestamp 1681620392
transform 1 0 736 0 1 770
box -8 -3 104 105
use INVX2  INVX2_287
timestamp 1681620392
transform -1 0 848 0 1 770
box -9 -3 26 105
use FILL  FILL_1097
timestamp 1681620392
transform 1 0 848 0 1 770
box -8 -3 16 105
use FILL  FILL_1098
timestamp 1681620392
transform 1 0 856 0 1 770
box -8 -3 16 105
use FILL  FILL_1099
timestamp 1681620392
transform 1 0 864 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_3779
timestamp 1681620392
transform 1 0 900 0 1 775
box -3 -3 3 3
use OAI21X1  OAI21X1_251
timestamp 1681620392
transform -1 0 904 0 1 770
box -8 -3 34 105
use INVX2  INVX2_288
timestamp 1681620392
transform -1 0 920 0 1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_238
timestamp 1681620392
transform -1 0 1016 0 1 770
box -8 -3 104 105
use FILL  FILL_1100
timestamp 1681620392
transform 1 0 1016 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_3780
timestamp 1681620392
transform 1 0 1052 0 1 775
box -3 -3 3 3
use AOI21X1  AOI21X1_28
timestamp 1681620392
transform -1 0 1056 0 1 770
box -7 -3 39 105
use FILL  FILL_1101
timestamp 1681620392
transform 1 0 1056 0 1 770
box -8 -3 16 105
use INVX2  INVX2_289
timestamp 1681620392
transform -1 0 1080 0 1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_239
timestamp 1681620392
transform -1 0 1176 0 1 770
box -8 -3 104 105
use M3_M2  M3_M2_3781
timestamp 1681620392
transform 1 0 1188 0 1 775
box -3 -3 3 3
use FILL  FILL_1102
timestamp 1681620392
transform 1 0 1176 0 1 770
box -8 -3 16 105
use FILL  FILL_1103
timestamp 1681620392
transform 1 0 1184 0 1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_253
timestamp 1681620392
transform 1 0 1192 0 1 770
box -8 -3 32 105
use OAI21X1  OAI21X1_252
timestamp 1681620392
transform 1 0 1216 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_253
timestamp 1681620392
transform 1 0 1248 0 1 770
box -8 -3 34 105
use NOR2X1  NOR2X1_83
timestamp 1681620392
transform 1 0 1280 0 1 770
box -8 -3 32 105
use FILL  FILL_1104
timestamp 1681620392
transform 1 0 1304 0 1 770
box -8 -3 16 105
use FILL  FILL_1105
timestamp 1681620392
transform 1 0 1312 0 1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_84
timestamp 1681620392
transform -1 0 1344 0 1 770
box -8 -3 32 105
use OAI21X1  OAI21X1_254
timestamp 1681620392
transform 1 0 1344 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_255
timestamp 1681620392
transform -1 0 1408 0 1 770
box -8 -3 34 105
use NAND2X1  NAND2X1_254
timestamp 1681620392
transform 1 0 1408 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_255
timestamp 1681620392
transform -1 0 1456 0 1 770
box -8 -3 32 105
use FILL  FILL_1106
timestamp 1681620392
transform 1 0 1456 0 1 770
box -8 -3 16 105
use INVX2  INVX2_290
timestamp 1681620392
transform -1 0 1480 0 1 770
box -9 -3 26 105
use OAI22X1  OAI22X1_82
timestamp 1681620392
transform 1 0 1480 0 1 770
box -8 -3 46 105
use M3_M2  M3_M2_3782
timestamp 1681620392
transform 1 0 1556 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_240
timestamp 1681620392
transform -1 0 1616 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_241
timestamp 1681620392
transform 1 0 1616 0 1 770
box -8 -3 104 105
use FILL  FILL_1107
timestamp 1681620392
transform 1 0 1712 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_3783
timestamp 1681620392
transform 1 0 1740 0 1 775
box -3 -3 3 3
use OAI22X1  OAI22X1_83
timestamp 1681620392
transform 1 0 1720 0 1 770
box -8 -3 46 105
use M3_M2  M3_M2_3784
timestamp 1681620392
transform 1 0 1772 0 1 775
box -3 -3 3 3
use NAND2X1  NAND2X1_256
timestamp 1681620392
transform -1 0 1784 0 1 770
box -8 -3 32 105
use INVX2  INVX2_291
timestamp 1681620392
transform 1 0 1784 0 1 770
box -9 -3 26 105
use M3_M2  M3_M2_3785
timestamp 1681620392
transform 1 0 1820 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3786
timestamp 1681620392
transform 1 0 1876 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_242
timestamp 1681620392
transform -1 0 1896 0 1 770
box -8 -3 104 105
use OAI21X1  OAI21X1_256
timestamp 1681620392
transform 1 0 1896 0 1 770
box -8 -3 34 105
use NAND2X1  NAND2X1_257
timestamp 1681620392
transform -1 0 1952 0 1 770
box -8 -3 32 105
use FILL  FILL_1108
timestamp 1681620392
transform 1 0 1952 0 1 770
box -8 -3 16 105
use FILL  FILL_1129
timestamp 1681620392
transform 1 0 1960 0 1 770
box -8 -3 16 105
use FILL  FILL_1131
timestamp 1681620392
transform 1 0 1968 0 1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_262
timestamp 1681620392
transform -1 0 2000 0 1 770
box -8 -3 32 105
use M3_M2  M3_M2_3787
timestamp 1681620392
transform 1 0 2100 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_249
timestamp 1681620392
transform 1 0 2000 0 1 770
box -8 -3 104 105
use FILL  FILL_1132
timestamp 1681620392
transform 1 0 2096 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_3788
timestamp 1681620392
transform 1 0 2116 0 1 775
box -3 -3 3 3
use OAI22X1  OAI22X1_87
timestamp 1681620392
transform -1 0 2144 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_88
timestamp 1681620392
transform -1 0 2184 0 1 770
box -8 -3 46 105
use INVX2  INVX2_297
timestamp 1681620392
transform 1 0 2184 0 1 770
box -9 -3 26 105
use OAI21X1  OAI21X1_258
timestamp 1681620392
transform 1 0 2200 0 1 770
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_250
timestamp 1681620392
transform 1 0 2232 0 1 770
box -8 -3 104 105
use FILL  FILL_1133
timestamp 1681620392
transform 1 0 2328 0 1 770
box -8 -3 16 105
use FILL  FILL_1134
timestamp 1681620392
transform 1 0 2336 0 1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_263
timestamp 1681620392
transform 1 0 2344 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_264
timestamp 1681620392
transform 1 0 2368 0 1 770
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_251
timestamp 1681620392
transform 1 0 2392 0 1 770
box -8 -3 104 105
use FILL  FILL_1135
timestamp 1681620392
transform 1 0 2488 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_259
timestamp 1681620392
transform -1 0 2528 0 1 770
box -8 -3 34 105
use FILL  FILL_1136
timestamp 1681620392
transform 1 0 2528 0 1 770
box -8 -3 16 105
use FILL  FILL_1137
timestamp 1681620392
transform 1 0 2536 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_260
timestamp 1681620392
transform -1 0 2576 0 1 770
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_252
timestamp 1681620392
transform 1 0 2576 0 1 770
box -8 -3 104 105
use INVX2  INVX2_298
timestamp 1681620392
transform -1 0 2688 0 1 770
box -9 -3 26 105
use FILL  FILL_1138
timestamp 1681620392
transform 1 0 2688 0 1 770
box -8 -3 16 105
use FILL  FILL_1139
timestamp 1681620392
transform 1 0 2696 0 1 770
box -8 -3 16 105
use FILL  FILL_1140
timestamp 1681620392
transform 1 0 2704 0 1 770
box -8 -3 16 105
use FILL  FILL_1141
timestamp 1681620392
transform 1 0 2712 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_264
timestamp 1681620392
transform 1 0 2720 0 1 770
box -8 -3 34 105
use FILL  FILL_1159
timestamp 1681620392
transform 1 0 2752 0 1 770
box -8 -3 16 105
use FILL  FILL_1160
timestamp 1681620392
transform 1 0 2760 0 1 770
box -8 -3 16 105
use FILL  FILL_1161
timestamp 1681620392
transform 1 0 2768 0 1 770
box -8 -3 16 105
use FILL  FILL_1162
timestamp 1681620392
transform 1 0 2776 0 1 770
box -8 -3 16 105
use FILL  FILL_1163
timestamp 1681620392
transform 1 0 2784 0 1 770
box -8 -3 16 105
use FILL  FILL_1164
timestamp 1681620392
transform 1 0 2792 0 1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_88
timestamp 1681620392
transform 1 0 2800 0 1 770
box -8 -3 32 105
use M3_M2  M3_M2_3789
timestamp 1681620392
transform 1 0 2836 0 1 775
box -3 -3 3 3
use FILL  FILL_1165
timestamp 1681620392
transform 1 0 2824 0 1 770
box -8 -3 16 105
use FILL  FILL_1166
timestamp 1681620392
transform 1 0 2832 0 1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_267
timestamp 1681620392
transform 1 0 2840 0 1 770
box -8 -3 32 105
use OAI21X1  OAI21X1_265
timestamp 1681620392
transform 1 0 2864 0 1 770
box -8 -3 34 105
use M3_M2  M3_M2_3790
timestamp 1681620392
transform 1 0 2916 0 1 775
box -3 -3 3 3
use INVX2  INVX2_302
timestamp 1681620392
transform 1 0 2896 0 1 770
box -9 -3 26 105
use NAND3X1  NAND3X1_96
timestamp 1681620392
transform 1 0 2912 0 1 770
box -8 -3 40 105
use M3_M2  M3_M2_3791
timestamp 1681620392
transform 1 0 2972 0 1 775
box -3 -3 3 3
use NOR2X1  NOR2X1_89
timestamp 1681620392
transform -1 0 2968 0 1 770
box -8 -3 32 105
use FILL  FILL_1170
timestamp 1681620392
transform 1 0 2968 0 1 770
box -8 -3 16 105
use FILL  FILL_1171
timestamp 1681620392
transform 1 0 2976 0 1 770
box -8 -3 16 105
use INVX2  INVX2_303
timestamp 1681620392
transform 1 0 2984 0 1 770
box -9 -3 26 105
use FILL  FILL_1172
timestamp 1681620392
transform 1 0 3000 0 1 770
box -8 -3 16 105
use FILL  FILL_1173
timestamp 1681620392
transform 1 0 3008 0 1 770
box -8 -3 16 105
use Project_Top_VIA0  Project_Top_VIA0_45
timestamp 1681620392
transform 1 0 3043 0 1 770
box -10 -3 10 3
use M2_M1  M2_M1_4360
timestamp 1681620392
transform 1 0 84 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3792
timestamp 1681620392
transform 1 0 220 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3793
timestamp 1681620392
transform 1 0 268 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_4361
timestamp 1681620392
transform 1 0 268 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4436
timestamp 1681620392
transform 1 0 132 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4437
timestamp 1681620392
transform 1 0 172 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4438
timestamp 1681620392
transform 1 0 180 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4439
timestamp 1681620392
transform 1 0 188 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4440
timestamp 1681620392
transform 1 0 244 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3874
timestamp 1681620392
transform 1 0 172 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3802
timestamp 1681620392
transform 1 0 300 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_4352
timestamp 1681620392
transform 1 0 316 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4362
timestamp 1681620392
transform 1 0 300 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3902
timestamp 1681620392
transform 1 0 292 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_4441
timestamp 1681620392
transform 1 0 316 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3803
timestamp 1681620392
transform 1 0 332 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_4353
timestamp 1681620392
transform 1 0 332 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4363
timestamp 1681620392
transform 1 0 340 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4442
timestamp 1681620392
transform 1 0 340 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3875
timestamp 1681620392
transform 1 0 340 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3903
timestamp 1681620392
transform 1 0 340 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_4354
timestamp 1681620392
transform 1 0 388 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4364
timestamp 1681620392
transform 1 0 364 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4365
timestamp 1681620392
transform 1 0 372 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4443
timestamp 1681620392
transform 1 0 356 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4444
timestamp 1681620392
transform 1 0 388 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4445
timestamp 1681620392
transform 1 0 396 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3876
timestamp 1681620392
transform 1 0 388 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_4366
timestamp 1681620392
transform 1 0 404 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4367
timestamp 1681620392
transform 1 0 452 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4446
timestamp 1681620392
transform 1 0 428 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4512
timestamp 1681620392
transform 1 0 420 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4530
timestamp 1681620392
transform 1 0 412 0 1 705
box -2 -2 2 2
use M3_M2  M3_M2_3913
timestamp 1681620392
transform 1 0 420 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_4513
timestamp 1681620392
transform 1 0 444 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3904
timestamp 1681620392
transform 1 0 444 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_4447
timestamp 1681620392
transform 1 0 468 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4368
timestamp 1681620392
transform 1 0 484 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4369
timestamp 1681620392
transform 1 0 516 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4448
timestamp 1681620392
transform 1 0 516 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4370
timestamp 1681620392
transform 1 0 532 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3857
timestamp 1681620392
transform 1 0 532 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_4449
timestamp 1681620392
transform 1 0 540 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4371
timestamp 1681620392
transform 1 0 556 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4514
timestamp 1681620392
transform 1 0 532 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3877
timestamp 1681620392
transform 1 0 548 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_4515
timestamp 1681620392
transform 1 0 556 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3914
timestamp 1681620392
transform 1 0 532 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_4372
timestamp 1681620392
transform 1 0 588 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4373
timestamp 1681620392
transform 1 0 596 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3858
timestamp 1681620392
transform 1 0 596 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_4450
timestamp 1681620392
transform 1 0 620 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4516
timestamp 1681620392
transform 1 0 596 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4517
timestamp 1681620392
transform 1 0 612 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3878
timestamp 1681620392
transform 1 0 620 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_4451
timestamp 1681620392
transform 1 0 636 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4518
timestamp 1681620392
transform 1 0 628 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4531
timestamp 1681620392
transform 1 0 620 0 1 705
box -2 -2 2 2
use M3_M2  M3_M2_3915
timestamp 1681620392
transform 1 0 628 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3822
timestamp 1681620392
transform 1 0 668 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_4374
timestamp 1681620392
transform 1 0 668 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4452
timestamp 1681620392
transform 1 0 660 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4519
timestamp 1681620392
transform 1 0 660 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3823
timestamp 1681620392
transform 1 0 708 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_4520
timestamp 1681620392
transform 1 0 700 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3794
timestamp 1681620392
transform 1 0 724 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3804
timestamp 1681620392
transform 1 0 724 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3795
timestamp 1681620392
transform 1 0 764 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3824
timestamp 1681620392
transform 1 0 748 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3825
timestamp 1681620392
transform 1 0 804 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_4375
timestamp 1681620392
transform 1 0 724 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4376
timestamp 1681620392
transform 1 0 732 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4377
timestamp 1681620392
transform 1 0 748 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4378
timestamp 1681620392
transform 1 0 764 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4379
timestamp 1681620392
transform 1 0 780 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4453
timestamp 1681620392
transform 1 0 740 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4454
timestamp 1681620392
transform 1 0 764 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4455
timestamp 1681620392
transform 1 0 804 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4456
timestamp 1681620392
transform 1 0 860 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4457
timestamp 1681620392
transform 1 0 868 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3879
timestamp 1681620392
transform 1 0 740 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3880
timestamp 1681620392
transform 1 0 764 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3905
timestamp 1681620392
transform 1 0 732 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3916
timestamp 1681620392
transform 1 0 748 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3881
timestamp 1681620392
transform 1 0 868 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3796
timestamp 1681620392
transform 1 0 892 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3805
timestamp 1681620392
transform 1 0 884 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_4355
timestamp 1681620392
transform 1 0 884 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4380
timestamp 1681620392
transform 1 0 876 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4381
timestamp 1681620392
transform 1 0 908 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4458
timestamp 1681620392
transform 1 0 884 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3859
timestamp 1681620392
transform 1 0 892 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_4459
timestamp 1681620392
transform 1 0 908 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4460
timestamp 1681620392
transform 1 0 916 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3882
timestamp 1681620392
transform 1 0 884 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3826
timestamp 1681620392
transform 1 0 924 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3827
timestamp 1681620392
transform 1 0 1020 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_4382
timestamp 1681620392
transform 1 0 924 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4383
timestamp 1681620392
transform 1 0 940 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3860
timestamp 1681620392
transform 1 0 924 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_4461
timestamp 1681620392
transform 1 0 964 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3861
timestamp 1681620392
transform 1 0 1012 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_4462
timestamp 1681620392
transform 1 0 1020 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3883
timestamp 1681620392
transform 1 0 964 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3797
timestamp 1681620392
transform 1 0 1052 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_4384
timestamp 1681620392
transform 1 0 1052 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4385
timestamp 1681620392
transform 1 0 1068 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4463
timestamp 1681620392
transform 1 0 1044 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4464
timestamp 1681620392
transform 1 0 1060 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3862
timestamp 1681620392
transform 1 0 1068 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3884
timestamp 1681620392
transform 1 0 1076 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_4386
timestamp 1681620392
transform 1 0 1100 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4465
timestamp 1681620392
transform 1 0 1092 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3845
timestamp 1681620392
transform 1 0 1108 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3863
timestamp 1681620392
transform 1 0 1124 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3828
timestamp 1681620392
transform 1 0 1148 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3806
timestamp 1681620392
transform 1 0 1172 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_4356
timestamp 1681620392
transform 1 0 1172 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4387
timestamp 1681620392
transform 1 0 1140 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3846
timestamp 1681620392
transform 1 0 1156 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_4388
timestamp 1681620392
transform 1 0 1164 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4466
timestamp 1681620392
transform 1 0 1132 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4467
timestamp 1681620392
transform 1 0 1148 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4521
timestamp 1681620392
transform 1 0 1124 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3885
timestamp 1681620392
transform 1 0 1132 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_4468
timestamp 1681620392
transform 1 0 1172 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3829
timestamp 1681620392
transform 1 0 1196 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_4389
timestamp 1681620392
transform 1 0 1196 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3807
timestamp 1681620392
transform 1 0 1220 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_4469
timestamp 1681620392
transform 1 0 1212 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4390
timestamp 1681620392
transform 1 0 1220 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3808
timestamp 1681620392
transform 1 0 1252 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3847
timestamp 1681620392
transform 1 0 1252 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3864
timestamp 1681620392
transform 1 0 1236 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_4470
timestamp 1681620392
transform 1 0 1252 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4471
timestamp 1681620392
transform 1 0 1260 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4522
timestamp 1681620392
transform 1 0 1252 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3906
timestamp 1681620392
transform 1 0 1244 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3809
timestamp 1681620392
transform 1 0 1292 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_4357
timestamp 1681620392
transform 1 0 1284 0 1 745
box -2 -2 2 2
use M3_M2  M3_M2_3848
timestamp 1681620392
transform 1 0 1284 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3810
timestamp 1681620392
transform 1 0 1332 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3811
timestamp 1681620392
transform 1 0 1396 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3830
timestamp 1681620392
transform 1 0 1308 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_4391
timestamp 1681620392
transform 1 0 1292 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4392
timestamp 1681620392
transform 1 0 1300 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3917
timestamp 1681620392
transform 1 0 1284 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_4393
timestamp 1681620392
transform 1 0 1396 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4472
timestamp 1681620392
transform 1 0 1308 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4473
timestamp 1681620392
transform 1 0 1372 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3921
timestamp 1681620392
transform 1 0 1388 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3922
timestamp 1681620392
transform 1 0 1420 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3798
timestamp 1681620392
transform 1 0 1524 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_4358
timestamp 1681620392
transform 1 0 1524 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4394
timestamp 1681620392
transform 1 0 1436 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4395
timestamp 1681620392
transform 1 0 1524 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4474
timestamp 1681620392
transform 1 0 1484 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4475
timestamp 1681620392
transform 1 0 1516 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3907
timestamp 1681620392
transform 1 0 1436 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3831
timestamp 1681620392
transform 1 0 1572 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_4359
timestamp 1681620392
transform 1 0 1580 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4396
timestamp 1681620392
transform 1 0 1564 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3849
timestamp 1681620392
transform 1 0 1572 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_4476
timestamp 1681620392
transform 1 0 1548 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4477
timestamp 1681620392
transform 1 0 1556 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3886
timestamp 1681620392
transform 1 0 1556 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3812
timestamp 1681620392
transform 1 0 1604 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_4478
timestamp 1681620392
transform 1 0 1596 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3887
timestamp 1681620392
transform 1 0 1596 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_4397
timestamp 1681620392
transform 1 0 1612 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4479
timestamp 1681620392
transform 1 0 1636 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3888
timestamp 1681620392
transform 1 0 1636 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3918
timestamp 1681620392
transform 1 0 1612 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3850
timestamp 1681620392
transform 1 0 1708 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_4398
timestamp 1681620392
transform 1 0 1716 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4480
timestamp 1681620392
transform 1 0 1708 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4481
timestamp 1681620392
transform 1 0 1732 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3889
timestamp 1681620392
transform 1 0 1732 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3813
timestamp 1681620392
transform 1 0 1756 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3814
timestamp 1681620392
transform 1 0 1844 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3832
timestamp 1681620392
transform 1 0 1756 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3833
timestamp 1681620392
transform 1 0 1804 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_4399
timestamp 1681620392
transform 1 0 1756 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4400
timestamp 1681620392
transform 1 0 1844 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4401
timestamp 1681620392
transform 1 0 1860 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3851
timestamp 1681620392
transform 1 0 1868 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3799
timestamp 1681620392
transform 1 0 1900 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_4402
timestamp 1681620392
transform 1 0 1876 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4403
timestamp 1681620392
transform 1 0 1884 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3865
timestamp 1681620392
transform 1 0 1756 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_4482
timestamp 1681620392
transform 1 0 1804 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4483
timestamp 1681620392
transform 1 0 1836 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3866
timestamp 1681620392
transform 1 0 1844 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_4484
timestamp 1681620392
transform 1 0 1852 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4485
timestamp 1681620392
transform 1 0 1868 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4486
timestamp 1681620392
transform 1 0 1876 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3890
timestamp 1681620392
transform 1 0 1876 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3908
timestamp 1681620392
transform 1 0 1884 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3834
timestamp 1681620392
transform 1 0 1908 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_4404
timestamp 1681620392
transform 1 0 1908 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4405
timestamp 1681620392
transform 1 0 1916 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3867
timestamp 1681620392
transform 1 0 1916 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3891
timestamp 1681620392
transform 1 0 1916 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3800
timestamp 1681620392
transform 1 0 1940 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_4406
timestamp 1681620392
transform 1 0 1948 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4523
timestamp 1681620392
transform 1 0 1932 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3923
timestamp 1681620392
transform 1 0 1892 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3892
timestamp 1681620392
transform 1 0 1940 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3909
timestamp 1681620392
transform 1 0 1940 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3852
timestamp 1681620392
transform 1 0 1980 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_4407
timestamp 1681620392
transform 1 0 1988 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4487
timestamp 1681620392
transform 1 0 1980 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4524
timestamp 1681620392
transform 1 0 2012 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3835
timestamp 1681620392
transform 1 0 2028 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3801
timestamp 1681620392
transform 1 0 2052 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3815
timestamp 1681620392
transform 1 0 2044 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_4408
timestamp 1681620392
transform 1 0 2036 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3836
timestamp 1681620392
transform 1 0 2084 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_4409
timestamp 1681620392
transform 1 0 2068 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4488
timestamp 1681620392
transform 1 0 2116 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3893
timestamp 1681620392
transform 1 0 2068 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3894
timestamp 1681620392
transform 1 0 2140 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3924
timestamp 1681620392
transform 1 0 2076 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3853
timestamp 1681620392
transform 1 0 2164 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_4489
timestamp 1681620392
transform 1 0 2172 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3895
timestamp 1681620392
transform 1 0 2172 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3854
timestamp 1681620392
transform 1 0 2220 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_4410
timestamp 1681620392
transform 1 0 2268 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4490
timestamp 1681620392
transform 1 0 2188 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4491
timestamp 1681620392
transform 1 0 2220 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4411
timestamp 1681620392
transform 1 0 2284 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4492
timestamp 1681620392
transform 1 0 2284 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3896
timestamp 1681620392
transform 1 0 2284 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3925
timestamp 1681620392
transform 1 0 2276 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_4412
timestamp 1681620392
transform 1 0 2324 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4525
timestamp 1681620392
transform 1 0 2332 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3926
timestamp 1681620392
transform 1 0 2308 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3927
timestamp 1681620392
transform 1 0 2332 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_4413
timestamp 1681620392
transform 1 0 2364 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4414
timestamp 1681620392
transform 1 0 2372 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4493
timestamp 1681620392
transform 1 0 2388 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3816
timestamp 1681620392
transform 1 0 2412 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_4415
timestamp 1681620392
transform 1 0 2412 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_3855
timestamp 1681620392
transform 1 0 2460 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3856
timestamp 1681620392
transform 1 0 2492 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3868
timestamp 1681620392
transform 1 0 2412 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_4494
timestamp 1681620392
transform 1 0 2460 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4526
timestamp 1681620392
transform 1 0 2396 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3910
timestamp 1681620392
transform 1 0 2452 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3837
timestamp 1681620392
transform 1 0 2516 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_4416
timestamp 1681620392
transform 1 0 2516 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4495
timestamp 1681620392
transform 1 0 2508 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3817
timestamp 1681620392
transform 1 0 2540 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3818
timestamp 1681620392
transform 1 0 2556 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3819
timestamp 1681620392
transform 1 0 2588 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3838
timestamp 1681620392
transform 1 0 2580 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_4417
timestamp 1681620392
transform 1 0 2540 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4418
timestamp 1681620392
transform 1 0 2556 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4496
timestamp 1681620392
transform 1 0 2532 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4527
timestamp 1681620392
transform 1 0 2516 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4497
timestamp 1681620392
transform 1 0 2580 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3897
timestamp 1681620392
transform 1 0 2540 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3911
timestamp 1681620392
transform 1 0 2532 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_4498
timestamp 1681620392
transform 1 0 2652 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4499
timestamp 1681620392
transform 1 0 2660 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3898
timestamp 1681620392
transform 1 0 2652 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3820
timestamp 1681620392
transform 1 0 2676 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3821
timestamp 1681620392
transform 1 0 2716 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3839
timestamp 1681620392
transform 1 0 2684 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3840
timestamp 1681620392
transform 1 0 2708 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_4419
timestamp 1681620392
transform 1 0 2676 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4420
timestamp 1681620392
transform 1 0 2692 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4421
timestamp 1681620392
transform 1 0 2708 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4422
timestamp 1681620392
transform 1 0 2716 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4500
timestamp 1681620392
transform 1 0 2700 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3869
timestamp 1681620392
transform 1 0 2708 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_4501
timestamp 1681620392
transform 1 0 2716 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3841
timestamp 1681620392
transform 1 0 2764 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3842
timestamp 1681620392
transform 1 0 2788 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_4423
timestamp 1681620392
transform 1 0 2740 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4424
timestamp 1681620392
transform 1 0 2756 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4425
timestamp 1681620392
transform 1 0 2764 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4426
timestamp 1681620392
transform 1 0 2780 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4427
timestamp 1681620392
transform 1 0 2796 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4428
timestamp 1681620392
transform 1 0 2804 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4502
timestamp 1681620392
transform 1 0 2748 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3870
timestamp 1681620392
transform 1 0 2756 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_4503
timestamp 1681620392
transform 1 0 2764 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4504
timestamp 1681620392
transform 1 0 2788 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3871
timestamp 1681620392
transform 1 0 2796 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3899
timestamp 1681620392
transform 1 0 2764 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3843
timestamp 1681620392
transform 1 0 2836 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_4429
timestamp 1681620392
transform 1 0 2836 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4505
timestamp 1681620392
transform 1 0 2812 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4506
timestamp 1681620392
transform 1 0 2828 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3900
timestamp 1681620392
transform 1 0 2828 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3919
timestamp 1681620392
transform 1 0 2812 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_4430
timestamp 1681620392
transform 1 0 2852 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4507
timestamp 1681620392
transform 1 0 2852 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3912
timestamp 1681620392
transform 1 0 2852 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3920
timestamp 1681620392
transform 1 0 2852 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_4431
timestamp 1681620392
transform 1 0 2868 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4508
timestamp 1681620392
transform 1 0 2876 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3872
timestamp 1681620392
transform 1 0 2884 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_4432
timestamp 1681620392
transform 1 0 2908 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4433
timestamp 1681620392
transform 1 0 2916 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4434
timestamp 1681620392
transform 1 0 2932 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4509
timestamp 1681620392
transform 1 0 2900 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4528
timestamp 1681620392
transform 1 0 2892 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3901
timestamp 1681620392
transform 1 0 2900 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_4510
timestamp 1681620392
transform 1 0 2940 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_3844
timestamp 1681620392
transform 1 0 2996 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_4435
timestamp 1681620392
transform 1 0 3004 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4511
timestamp 1681620392
transform 1 0 2996 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4529
timestamp 1681620392
transform 1 0 2980 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_3873
timestamp 1681620392
transform 1 0 3004 0 1 725
box -3 -3 3 3
use Project_Top_VIA0  Project_Top_VIA0_46
timestamp 1681620392
transform 1 0 24 0 1 670
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_235
timestamp 1681620392
transform 1 0 72 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_281
timestamp 1681620392
transform 1 0 168 0 -1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_236
timestamp 1681620392
transform -1 0 280 0 -1 770
box -8 -3 104 105
use FILL  FILL_1080
timestamp 1681620392
transform 1 0 280 0 -1 770
box -8 -3 16 105
use FILL  FILL_1081
timestamp 1681620392
transform 1 0 288 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_282
timestamp 1681620392
transform 1 0 296 0 -1 770
box -9 -3 26 105
use NOR2X1  NOR2X1_81
timestamp 1681620392
transform 1 0 312 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_82
timestamp 1681620392
transform 1 0 336 0 -1 770
box -8 -3 32 105
use AOI21X1  AOI21X1_27
timestamp 1681620392
transform 1 0 360 0 -1 770
box -7 -3 39 105
use INVX2  INVX2_283
timestamp 1681620392
transform -1 0 408 0 -1 770
box -9 -3 26 105
use FILL  FILL_1082
timestamp 1681620392
transform 1 0 408 0 -1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_93
timestamp 1681620392
transform 1 0 416 0 -1 770
box -8 -3 40 105
use INVX2  INVX2_284
timestamp 1681620392
transform 1 0 448 0 -1 770
box -9 -3 26 105
use FILL  FILL_1083
timestamp 1681620392
transform 1 0 464 0 -1 770
box -8 -3 16 105
use FILL  FILL_1084
timestamp 1681620392
transform 1 0 472 0 -1 770
box -8 -3 16 105
use FILL  FILL_1086
timestamp 1681620392
transform 1 0 480 0 -1 770
box -8 -3 16 105
use FILL  FILL_1093
timestamp 1681620392
transform 1 0 488 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_286
timestamp 1681620392
transform 1 0 496 0 -1 770
box -9 -3 26 105
use NAND2X1  NAND2X1_250
timestamp 1681620392
transform 1 0 512 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_251
timestamp 1681620392
transform 1 0 536 0 -1 770
box -8 -3 32 105
use OAI21X1  OAI21X1_248
timestamp 1681620392
transform 1 0 560 0 -1 770
box -8 -3 34 105
use NAND2X1  NAND2X1_252
timestamp 1681620392
transform 1 0 592 0 -1 770
box -8 -3 32 105
use FILL  FILL_1094
timestamp 1681620392
transform 1 0 616 0 -1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_95
timestamp 1681620392
transform 1 0 624 0 -1 770
box -8 -3 40 105
use FILL  FILL_1095
timestamp 1681620392
transform 1 0 656 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_249
timestamp 1681620392
transform 1 0 664 0 -1 770
box -8 -3 34 105
use FILL  FILL_1096
timestamp 1681620392
transform 1 0 696 0 -1 770
box -8 -3 16 105
use FILL  FILL_1109
timestamp 1681620392
transform 1 0 704 0 -1 770
box -8 -3 16 105
use FILL  FILL_1110
timestamp 1681620392
transform 1 0 712 0 -1 770
box -8 -3 16 105
use FILL  FILL_1111
timestamp 1681620392
transform 1 0 720 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_84
timestamp 1681620392
transform -1 0 768 0 -1 770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_243
timestamp 1681620392
transform 1 0 768 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_292
timestamp 1681620392
transform -1 0 880 0 -1 770
box -9 -3 26 105
use AOI21X1  AOI21X1_29
timestamp 1681620392
transform -1 0 912 0 -1 770
box -7 -3 39 105
use INVX2  INVX2_293
timestamp 1681620392
transform -1 0 928 0 -1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_244
timestamp 1681620392
transform 1 0 928 0 -1 770
box -8 -3 104 105
use FILL  FILL_1112
timestamp 1681620392
transform 1 0 1024 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_85
timestamp 1681620392
transform 1 0 1032 0 -1 770
box -8 -3 46 105
use FILL  FILL_1113
timestamp 1681620392
transform 1 0 1072 0 -1 770
box -8 -3 16 105
use FILL  FILL_1114
timestamp 1681620392
transform 1 0 1080 0 -1 770
box -8 -3 16 105
use FILL  FILL_1115
timestamp 1681620392
transform 1 0 1088 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_258
timestamp 1681620392
transform 1 0 1096 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_259
timestamp 1681620392
transform -1 0 1144 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_85
timestamp 1681620392
transform -1 0 1168 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_86
timestamp 1681620392
transform -1 0 1192 0 -1 770
box -8 -3 32 105
use INVX2  INVX2_294
timestamp 1681620392
transform 1 0 1192 0 -1 770
box -9 -3 26 105
use FILL  FILL_1116
timestamp 1681620392
transform 1 0 1208 0 -1 770
box -8 -3 16 105
use FILL  FILL_1117
timestamp 1681620392
transform 1 0 1216 0 -1 770
box -8 -3 16 105
use FILL  FILL_1118
timestamp 1681620392
transform 1 0 1224 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_260
timestamp 1681620392
transform 1 0 1232 0 -1 770
box -8 -3 32 105
use BUFX2  BUFX2_37
timestamp 1681620392
transform 1 0 1256 0 -1 770
box -5 -3 28 105
use FILL  FILL_1119
timestamp 1681620392
transform 1 0 1280 0 -1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_87
timestamp 1681620392
transform 1 0 1288 0 -1 770
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_245
timestamp 1681620392
transform -1 0 1408 0 -1 770
box -8 -3 104 105
use FILL  FILL_1120
timestamp 1681620392
transform 1 0 1408 0 -1 770
box -8 -3 16 105
use FILL  FILL_1121
timestamp 1681620392
transform 1 0 1416 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_246
timestamp 1681620392
transform 1 0 1424 0 -1 770
box -8 -3 104 105
use AOI21X1  AOI21X1_30
timestamp 1681620392
transform -1 0 1552 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_31
timestamp 1681620392
transform 1 0 1552 0 -1 770
box -7 -3 39 105
use FILL  FILL_1122
timestamp 1681620392
transform 1 0 1584 0 -1 770
box -8 -3 16 105
use FILL  FILL_1123
timestamp 1681620392
transform 1 0 1592 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_247
timestamp 1681620392
transform 1 0 1600 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_295
timestamp 1681620392
transform 1 0 1696 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_296
timestamp 1681620392
transform 1 0 1712 0 -1 770
box -9 -3 26 105
use FILL  FILL_1124
timestamp 1681620392
transform 1 0 1728 0 -1 770
box -8 -3 16 105
use FILL  FILL_1125
timestamp 1681620392
transform 1 0 1736 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_248
timestamp 1681620392
transform 1 0 1744 0 -1 770
box -8 -3 104 105
use OAI22X1  OAI22X1_86
timestamp 1681620392
transform -1 0 1880 0 -1 770
box -8 -3 46 105
use OAI21X1  OAI21X1_257
timestamp 1681620392
transform 1 0 1880 0 -1 770
box -8 -3 34 105
use NAND2X1  NAND2X1_261
timestamp 1681620392
transform 1 0 1912 0 -1 770
box -8 -3 32 105
use FILL  FILL_1126
timestamp 1681620392
transform 1 0 1936 0 -1 770
box -8 -3 16 105
use FILL  FILL_1127
timestamp 1681620392
transform 1 0 1944 0 -1 770
box -8 -3 16 105
use FILL  FILL_1128
timestamp 1681620392
transform 1 0 1952 0 -1 770
box -8 -3 16 105
use FILL  FILL_1130
timestamp 1681620392
transform 1 0 1960 0 -1 770
box -8 -3 16 105
use FILL  FILL_1142
timestamp 1681620392
transform 1 0 1968 0 -1 770
box -8 -3 16 105
use FILL  FILL_1143
timestamp 1681620392
transform 1 0 1976 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_261
timestamp 1681620392
transform 1 0 1984 0 -1 770
box -8 -3 34 105
use FILL  FILL_1144
timestamp 1681620392
transform 1 0 2016 0 -1 770
box -8 -3 16 105
use FILL  FILL_1145
timestamp 1681620392
transform 1 0 2024 0 -1 770
box -8 -3 16 105
use FILL  FILL_1146
timestamp 1681620392
transform 1 0 2032 0 -1 770
box -8 -3 16 105
use FILL  FILL_1147
timestamp 1681620392
transform 1 0 2040 0 -1 770
box -8 -3 16 105
use FILL  FILL_1148
timestamp 1681620392
transform 1 0 2048 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_253
timestamp 1681620392
transform 1 0 2056 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_299
timestamp 1681620392
transform 1 0 2152 0 -1 770
box -9 -3 26 105
use FILL  FILL_1149
timestamp 1681620392
transform 1 0 2168 0 -1 770
box -8 -3 16 105
use FILL  FILL_1150
timestamp 1681620392
transform 1 0 2176 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_254
timestamp 1681620392
transform -1 0 2280 0 -1 770
box -8 -3 104 105
use FILL  FILL_1151
timestamp 1681620392
transform 1 0 2280 0 -1 770
box -8 -3 16 105
use FILL  FILL_1152
timestamp 1681620392
transform 1 0 2288 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_262
timestamp 1681620392
transform 1 0 2296 0 -1 770
box -8 -3 34 105
use NAND2X1  NAND2X1_265
timestamp 1681620392
transform -1 0 2352 0 -1 770
box -8 -3 32 105
use FILL  FILL_1153
timestamp 1681620392
transform 1 0 2352 0 -1 770
box -8 -3 16 105
use FILL  FILL_1154
timestamp 1681620392
transform 1 0 2360 0 -1 770
box -8 -3 16 105
use FILL  FILL_1155
timestamp 1681620392
transform 1 0 2368 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_266
timestamp 1681620392
transform 1 0 2376 0 -1 770
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_255
timestamp 1681620392
transform 1 0 2400 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_300
timestamp 1681620392
transform 1 0 2496 0 -1 770
box -9 -3 26 105
use OAI21X1  OAI21X1_263
timestamp 1681620392
transform -1 0 2544 0 -1 770
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_256
timestamp 1681620392
transform 1 0 2544 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_301
timestamp 1681620392
transform 1 0 2640 0 -1 770
box -9 -3 26 105
use FILL  FILL_1156
timestamp 1681620392
transform 1 0 2656 0 -1 770
box -8 -3 16 105
use FILL  FILL_1157
timestamp 1681620392
transform 1 0 2664 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_89
timestamp 1681620392
transform 1 0 2672 0 -1 770
box -8 -3 46 105
use FILL  FILL_1158
timestamp 1681620392
transform 1 0 2712 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_90
timestamp 1681620392
transform 1 0 2720 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_91
timestamp 1681620392
transform 1 0 2760 0 -1 770
box -8 -3 46 105
use FILL  FILL_1167
timestamp 1681620392
transform 1 0 2800 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_42
timestamp 1681620392
transform -1 0 2848 0 -1 770
box -8 -3 46 105
use FILL  FILL_1168
timestamp 1681620392
transform 1 0 2848 0 -1 770
box -8 -3 16 105
use FILL  FILL_1169
timestamp 1681620392
transform 1 0 2856 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_266
timestamp 1681620392
transform 1 0 2864 0 -1 770
box -8 -3 34 105
use FILL  FILL_1174
timestamp 1681620392
transform 1 0 2896 0 -1 770
box -8 -3 16 105
use FILL  FILL_1175
timestamp 1681620392
transform 1 0 2904 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_92
timestamp 1681620392
transform 1 0 2912 0 -1 770
box -8 -3 46 105
use FILL  FILL_1176
timestamp 1681620392
transform 1 0 2952 0 -1 770
box -8 -3 16 105
use FILL  FILL_1177
timestamp 1681620392
transform 1 0 2960 0 -1 770
box -8 -3 16 105
use FILL  FILL_1178
timestamp 1681620392
transform 1 0 2968 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_267
timestamp 1681620392
transform -1 0 3008 0 -1 770
box -8 -3 34 105
use FILL  FILL_1179
timestamp 1681620392
transform 1 0 3008 0 -1 770
box -8 -3 16 105
use Project_Top_VIA0  Project_Top_VIA0_47
timestamp 1681620392
transform 1 0 3067 0 1 670
box -10 -3 10 3
use M3_M2  M3_M2_3965
timestamp 1681620392
transform 1 0 180 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4555
timestamp 1681620392
transform 1 0 140 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4556
timestamp 1681620392
transform 1 0 180 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4557
timestamp 1681620392
transform 1 0 188 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4640
timestamp 1681620392
transform 1 0 92 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4063
timestamp 1681620392
transform 1 0 164 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4015
timestamp 1681620392
transform 1 0 188 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_4724
timestamp 1681620392
transform 1 0 196 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_3966
timestamp 1681620392
transform 1 0 236 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3995
timestamp 1681620392
transform 1 0 228 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_4558
timestamp 1681620392
transform 1 0 236 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4641
timestamp 1681620392
transform 1 0 228 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4642
timestamp 1681620392
transform 1 0 236 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4725
timestamp 1681620392
transform 1 0 220 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_4030
timestamp 1681620392
transform 1 0 236 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4064
timestamp 1681620392
transform 1 0 244 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3967
timestamp 1681620392
transform 1 0 276 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4559
timestamp 1681620392
transform 1 0 268 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3968
timestamp 1681620392
transform 1 0 300 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4560
timestamp 1681620392
transform 1 0 284 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3996
timestamp 1681620392
transform 1 0 292 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_4561
timestamp 1681620392
transform 1 0 300 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_4031
timestamp 1681620392
transform 1 0 284 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4016
timestamp 1681620392
transform 1 0 300 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_4726
timestamp 1681620392
transform 1 0 300 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_3997
timestamp 1681620392
transform 1 0 316 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_4643
timestamp 1681620392
transform 1 0 316 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4017
timestamp 1681620392
transform 1 0 324 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3948
timestamp 1681620392
transform 1 0 348 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_4562
timestamp 1681620392
transform 1 0 348 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4644
timestamp 1681620392
transform 1 0 332 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4534
timestamp 1681620392
transform 1 0 380 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_3998
timestamp 1681620392
transform 1 0 380 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_4535
timestamp 1681620392
transform 1 0 396 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_3999
timestamp 1681620392
transform 1 0 396 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_4563
timestamp 1681620392
transform 1 0 404 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4645
timestamp 1681620392
transform 1 0 404 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4032
timestamp 1681620392
transform 1 0 404 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_4532
timestamp 1681620392
transform 1 0 420 0 1 635
box -2 -2 2 2
use M3_M2  M3_M2_3930
timestamp 1681620392
transform 1 0 484 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_4536
timestamp 1681620392
transform 1 0 436 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4537
timestamp 1681620392
transform 1 0 452 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4538
timestamp 1681620392
transform 1 0 476 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4564
timestamp 1681620392
transform 1 0 420 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_4000
timestamp 1681620392
transform 1 0 428 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_4565
timestamp 1681620392
transform 1 0 436 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4646
timestamp 1681620392
transform 1 0 420 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4001
timestamp 1681620392
transform 1 0 460 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3969
timestamp 1681620392
transform 1 0 492 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4566
timestamp 1681620392
transform 1 0 476 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4567
timestamp 1681620392
transform 1 0 484 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4568
timestamp 1681620392
transform 1 0 500 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4647
timestamp 1681620392
transform 1 0 460 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4018
timestamp 1681620392
transform 1 0 476 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_4065
timestamp 1681620392
transform 1 0 452 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_4648
timestamp 1681620392
transform 1 0 492 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4033
timestamp 1681620392
transform 1 0 500 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4019
timestamp 1681620392
transform 1 0 524 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_4727
timestamp 1681620392
transform 1 0 524 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_3949
timestamp 1681620392
transform 1 0 572 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_4539
timestamp 1681620392
transform 1 0 572 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4569
timestamp 1681620392
transform 1 0 572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4649
timestamp 1681620392
transform 1 0 556 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4034
timestamp 1681620392
transform 1 0 572 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_4650
timestamp 1681620392
transform 1 0 588 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4651
timestamp 1681620392
transform 1 0 596 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3931
timestamp 1681620392
transform 1 0 636 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3950
timestamp 1681620392
transform 1 0 620 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4020
timestamp 1681620392
transform 1 0 628 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3951
timestamp 1681620392
transform 1 0 660 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3952
timestamp 1681620392
transform 1 0 684 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_4540
timestamp 1681620392
transform 1 0 644 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4541
timestamp 1681620392
transform 1 0 660 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_3970
timestamp 1681620392
transform 1 0 668 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4002
timestamp 1681620392
transform 1 0 660 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_4542
timestamp 1681620392
transform 1 0 692 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4570
timestamp 1681620392
transform 1 0 668 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4571
timestamp 1681620392
transform 1 0 676 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4652
timestamp 1681620392
transform 1 0 636 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4653
timestamp 1681620392
transform 1 0 644 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4654
timestamp 1681620392
transform 1 0 660 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4035
timestamp 1681620392
transform 1 0 660 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4003
timestamp 1681620392
transform 1 0 692 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3971
timestamp 1681620392
transform 1 0 724 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4572
timestamp 1681620392
transform 1 0 700 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4573
timestamp 1681620392
transform 1 0 708 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4574
timestamp 1681620392
transform 1 0 724 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4655
timestamp 1681620392
transform 1 0 700 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4656
timestamp 1681620392
transform 1 0 716 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4657
timestamp 1681620392
transform 1 0 732 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4658
timestamp 1681620392
transform 1 0 748 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4036
timestamp 1681620392
transform 1 0 732 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4066
timestamp 1681620392
transform 1 0 716 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3972
timestamp 1681620392
transform 1 0 772 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4575
timestamp 1681620392
transform 1 0 772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4659
timestamp 1681620392
transform 1 0 772 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3973
timestamp 1681620392
transform 1 0 876 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4576
timestamp 1681620392
transform 1 0 812 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_4004
timestamp 1681620392
transform 1 0 860 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_4577
timestamp 1681620392
transform 1 0 868 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4578
timestamp 1681620392
transform 1 0 876 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4660
timestamp 1681620392
transform 1 0 788 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4037
timestamp 1681620392
transform 1 0 812 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_4543
timestamp 1681620392
transform 1 0 892 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_4005
timestamp 1681620392
transform 1 0 900 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4021
timestamp 1681620392
transform 1 0 892 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_4661
timestamp 1681620392
transform 1 0 900 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3953
timestamp 1681620392
transform 1 0 948 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3974
timestamp 1681620392
transform 1 0 932 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3975
timestamp 1681620392
transform 1 0 1036 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3976
timestamp 1681620392
transform 1 0 1060 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4579
timestamp 1681620392
transform 1 0 932 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4580
timestamp 1681620392
transform 1 0 972 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4581
timestamp 1681620392
transform 1 0 1028 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4582
timestamp 1681620392
transform 1 0 1036 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4583
timestamp 1681620392
transform 1 0 1044 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4662
timestamp 1681620392
transform 1 0 908 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4022
timestamp 1681620392
transform 1 0 916 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_4663
timestamp 1681620392
transform 1 0 932 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4664
timestamp 1681620392
transform 1 0 948 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4023
timestamp 1681620392
transform 1 0 972 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_4067
timestamp 1681620392
transform 1 0 932 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4006
timestamp 1681620392
transform 1 0 1052 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_4584
timestamp 1681620392
transform 1 0 1060 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_4007
timestamp 1681620392
transform 1 0 1068 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_4585
timestamp 1681620392
transform 1 0 1076 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3977
timestamp 1681620392
transform 1 0 1092 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4586
timestamp 1681620392
transform 1 0 1092 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4665
timestamp 1681620392
transform 1 0 1044 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4666
timestamp 1681620392
transform 1 0 1052 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4667
timestamp 1681620392
transform 1 0 1068 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4668
timestamp 1681620392
transform 1 0 1084 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4669
timestamp 1681620392
transform 1 0 1092 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4038
timestamp 1681620392
transform 1 0 1028 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4039
timestamp 1681620392
transform 1 0 1044 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3954
timestamp 1681620392
transform 1 0 1220 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3955
timestamp 1681620392
transform 1 0 1236 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_4587
timestamp 1681620392
transform 1 0 1124 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4588
timestamp 1681620392
transform 1 0 1140 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4589
timestamp 1681620392
transform 1 0 1172 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_4024
timestamp 1681620392
transform 1 0 1108 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_4670
timestamp 1681620392
transform 1 0 1116 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4671
timestamp 1681620392
transform 1 0 1132 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4040
timestamp 1681620392
transform 1 0 1092 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4041
timestamp 1681620392
transform 1 0 1116 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4068
timestamp 1681620392
transform 1 0 1124 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4025
timestamp 1681620392
transform 1 0 1172 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_4672
timestamp 1681620392
transform 1 0 1220 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4673
timestamp 1681620392
transform 1 0 1236 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4042
timestamp 1681620392
transform 1 0 1220 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4069
timestamp 1681620392
transform 1 0 1180 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_4590
timestamp 1681620392
transform 1 0 1252 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_4043
timestamp 1681620392
transform 1 0 1252 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3932
timestamp 1681620392
transform 1 0 1316 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3978
timestamp 1681620392
transform 1 0 1292 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4591
timestamp 1681620392
transform 1 0 1292 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4592
timestamp 1681620392
transform 1 0 1316 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4674
timestamp 1681620392
transform 1 0 1284 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4675
timestamp 1681620392
transform 1 0 1308 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4676
timestamp 1681620392
transform 1 0 1324 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4728
timestamp 1681620392
transform 1 0 1292 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_4044
timestamp 1681620392
transform 1 0 1316 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3956
timestamp 1681620392
transform 1 0 1340 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_4544
timestamp 1681620392
transform 1 0 1340 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4593
timestamp 1681620392
transform 1 0 1348 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4677
timestamp 1681620392
transform 1 0 1340 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4045
timestamp 1681620392
transform 1 0 1340 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3933
timestamp 1681620392
transform 1 0 1364 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3979
timestamp 1681620392
transform 1 0 1356 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3980
timestamp 1681620392
transform 1 0 1372 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3981
timestamp 1681620392
transform 1 0 1396 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4594
timestamp 1681620392
transform 1 0 1356 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4595
timestamp 1681620392
transform 1 0 1364 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3934
timestamp 1681620392
transform 1 0 1460 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_4545
timestamp 1681620392
transform 1 0 1468 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4596
timestamp 1681620392
transform 1 0 1388 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4597
timestamp 1681620392
transform 1 0 1396 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4598
timestamp 1681620392
transform 1 0 1420 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4599
timestamp 1681620392
transform 1 0 1436 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4600
timestamp 1681620392
transform 1 0 1460 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4601
timestamp 1681620392
transform 1 0 1484 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4678
timestamp 1681620392
transform 1 0 1372 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4679
timestamp 1681620392
transform 1 0 1396 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4680
timestamp 1681620392
transform 1 0 1412 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4681
timestamp 1681620392
transform 1 0 1428 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4682
timestamp 1681620392
transform 1 0 1460 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4683
timestamp 1681620392
transform 1 0 1468 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4729
timestamp 1681620392
transform 1 0 1388 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_4684
timestamp 1681620392
transform 1 0 1492 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4730
timestamp 1681620392
transform 1 0 1436 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_4046
timestamp 1681620392
transform 1 0 1460 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4047
timestamp 1681620392
transform 1 0 1484 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4070
timestamp 1681620392
transform 1 0 1436 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4071
timestamp 1681620392
transform 1 0 1492 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3935
timestamp 1681620392
transform 1 0 1540 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3982
timestamp 1681620392
transform 1 0 1532 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4602
timestamp 1681620392
transform 1 0 1516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4685
timestamp 1681620392
transform 1 0 1508 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4026
timestamp 1681620392
transform 1 0 1516 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_4603
timestamp 1681620392
transform 1 0 1540 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4686
timestamp 1681620392
transform 1 0 1532 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4731
timestamp 1681620392
transform 1 0 1516 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_3983
timestamp 1681620392
transform 1 0 1580 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4604
timestamp 1681620392
transform 1 0 1572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4605
timestamp 1681620392
transform 1 0 1580 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4687
timestamp 1681620392
transform 1 0 1556 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4027
timestamp 1681620392
transform 1 0 1572 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_4688
timestamp 1681620392
transform 1 0 1580 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4732
timestamp 1681620392
transform 1 0 1572 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_4072
timestamp 1681620392
transform 1 0 1580 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_4546
timestamp 1681620392
transform 1 0 1604 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4606
timestamp 1681620392
transform 1 0 1644 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4689
timestamp 1681620392
transform 1 0 1604 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4690
timestamp 1681620392
transform 1 0 1620 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4048
timestamp 1681620392
transform 1 0 1604 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4049
timestamp 1681620392
transform 1 0 1644 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3984
timestamp 1681620392
transform 1 0 1716 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4607
timestamp 1681620392
transform 1 0 1708 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4608
timestamp 1681620392
transform 1 0 1716 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4691
timestamp 1681620392
transform 1 0 1724 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4692
timestamp 1681620392
transform 1 0 1740 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3985
timestamp 1681620392
transform 1 0 1788 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4609
timestamp 1681620392
transform 1 0 1756 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4610
timestamp 1681620392
transform 1 0 1772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4611
timestamp 1681620392
transform 1 0 1780 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4693
timestamp 1681620392
transform 1 0 1764 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4050
timestamp 1681620392
transform 1 0 1764 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4073
timestamp 1681620392
transform 1 0 1756 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_4694
timestamp 1681620392
transform 1 0 1788 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4008
timestamp 1681620392
transform 1 0 1804 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_4612
timestamp 1681620392
transform 1 0 1828 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_4009
timestamp 1681620392
transform 1 0 1844 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_4695
timestamp 1681620392
transform 1 0 1804 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4051
timestamp 1681620392
transform 1 0 1828 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4074
timestamp 1681620392
transform 1 0 1804 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3928
timestamp 1681620392
transform 1 0 1900 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3986
timestamp 1681620392
transform 1 0 1908 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3929
timestamp 1681620392
transform 1 0 1948 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3941
timestamp 1681620392
transform 1 0 1948 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3957
timestamp 1681620392
transform 1 0 1940 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_4547
timestamp 1681620392
transform 1 0 1940 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4548
timestamp 1681620392
transform 1 0 1948 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4613
timestamp 1681620392
transform 1 0 1908 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4614
timestamp 1681620392
transform 1 0 1924 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4615
timestamp 1681620392
transform 1 0 1940 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4696
timestamp 1681620392
transform 1 0 1916 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4010
timestamp 1681620392
transform 1 0 1956 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3942
timestamp 1681620392
transform 1 0 2084 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3958
timestamp 1681620392
transform 1 0 2068 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4011
timestamp 1681620392
transform 1 0 1980 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_4616
timestamp 1681620392
transform 1 0 2004 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4617
timestamp 1681620392
transform 1 0 2060 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4618
timestamp 1681620392
transform 1 0 2068 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4697
timestamp 1681620392
transform 1 0 1948 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4698
timestamp 1681620392
transform 1 0 1964 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4699
timestamp 1681620392
transform 1 0 1980 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4052
timestamp 1681620392
transform 1 0 1948 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4028
timestamp 1681620392
transform 1 0 2020 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_4700
timestamp 1681620392
transform 1 0 2068 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4053
timestamp 1681620392
transform 1 0 2004 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4075
timestamp 1681620392
transform 1 0 2068 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_4549
timestamp 1681620392
transform 1 0 2084 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_4012
timestamp 1681620392
transform 1 0 2092 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3943
timestamp 1681620392
transform 1 0 2204 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3987
timestamp 1681620392
transform 1 0 2124 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4619
timestamp 1681620392
transform 1 0 2100 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4620
timestamp 1681620392
transform 1 0 2124 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4621
timestamp 1681620392
transform 1 0 2164 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4701
timestamp 1681620392
transform 1 0 2092 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4029
timestamp 1681620392
transform 1 0 2100 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_4702
timestamp 1681620392
transform 1 0 2108 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4703
timestamp 1681620392
transform 1 0 2124 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4704
timestamp 1681620392
transform 1 0 2140 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4054
timestamp 1681620392
transform 1 0 2108 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4055
timestamp 1681620392
transform 1 0 2164 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3988
timestamp 1681620392
transform 1 0 2236 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4622
timestamp 1681620392
transform 1 0 2236 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4705
timestamp 1681620392
transform 1 0 2244 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4550
timestamp 1681620392
transform 1 0 2276 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_3936
timestamp 1681620392
transform 1 0 2364 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3937
timestamp 1681620392
transform 1 0 2388 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_4623
timestamp 1681620392
transform 1 0 2332 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4624
timestamp 1681620392
transform 1 0 2388 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4706
timestamp 1681620392
transform 1 0 2276 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4707
timestamp 1681620392
transform 1 0 2292 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4708
timestamp 1681620392
transform 1 0 2308 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4709
timestamp 1681620392
transform 1 0 2396 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4056
timestamp 1681620392
transform 1 0 2292 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4057
timestamp 1681620392
transform 1 0 2372 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4076
timestamp 1681620392
transform 1 0 2396 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_4533
timestamp 1681620392
transform 1 0 2420 0 1 635
box -2 -2 2 2
use M3_M2  M3_M2_3989
timestamp 1681620392
transform 1 0 2420 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4625
timestamp 1681620392
transform 1 0 2420 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4710
timestamp 1681620392
transform 1 0 2412 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4058
timestamp 1681620392
transform 1 0 2420 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3944
timestamp 1681620392
transform 1 0 2436 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3959
timestamp 1681620392
transform 1 0 2444 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_4551
timestamp 1681620392
transform 1 0 2436 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_4013
timestamp 1681620392
transform 1 0 2436 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_4626
timestamp 1681620392
transform 1 0 2444 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4711
timestamp 1681620392
transform 1 0 2436 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4077
timestamp 1681620392
transform 1 0 2412 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4078
timestamp 1681620392
transform 1 0 2428 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3945
timestamp 1681620392
transform 1 0 2460 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_4552
timestamp 1681620392
transform 1 0 2460 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_3938
timestamp 1681620392
transform 1 0 2492 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3946
timestamp 1681620392
transform 1 0 2484 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_4627
timestamp 1681620392
transform 1 0 2484 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4628
timestamp 1681620392
transform 1 0 2492 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_3960
timestamp 1681620392
transform 1 0 2508 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_4553
timestamp 1681620392
transform 1 0 2508 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_3990
timestamp 1681620392
transform 1 0 2516 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4059
timestamp 1681620392
transform 1 0 2524 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_4712
timestamp 1681620392
transform 1 0 2540 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4629
timestamp 1681620392
transform 1 0 2564 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4713
timestamp 1681620392
transform 1 0 2548 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3947
timestamp 1681620392
transform 1 0 2636 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_4554
timestamp 1681620392
transform 1 0 2636 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_3991
timestamp 1681620392
transform 1 0 2668 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4630
timestamp 1681620392
transform 1 0 2660 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4714
timestamp 1681620392
transform 1 0 2660 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3961
timestamp 1681620392
transform 1 0 2692 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_4631
timestamp 1681620392
transform 1 0 2692 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4632
timestamp 1681620392
transform 1 0 2700 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4715
timestamp 1681620392
transform 1 0 2676 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4060
timestamp 1681620392
transform 1 0 2676 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3939
timestamp 1681620392
transform 1 0 2716 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3962
timestamp 1681620392
transform 1 0 2724 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3992
timestamp 1681620392
transform 1 0 2724 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4716
timestamp 1681620392
transform 1 0 2732 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4633
timestamp 1681620392
transform 1 0 2772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4717
timestamp 1681620392
transform 1 0 2820 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4061
timestamp 1681620392
transform 1 0 2772 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3940
timestamp 1681620392
transform 1 0 2844 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3993
timestamp 1681620392
transform 1 0 2868 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4634
timestamp 1681620392
transform 1 0 2852 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4718
timestamp 1681620392
transform 1 0 2844 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4014
timestamp 1681620392
transform 1 0 2860 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3963
timestamp 1681620392
transform 1 0 2892 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_4635
timestamp 1681620392
transform 1 0 2868 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4636
timestamp 1681620392
transform 1 0 2884 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4719
timestamp 1681620392
transform 1 0 2860 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4720
timestamp 1681620392
transform 1 0 2876 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_3964
timestamp 1681620392
transform 1 0 2940 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3994
timestamp 1681620392
transform 1 0 2932 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_4637
timestamp 1681620392
transform 1 0 2916 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4638
timestamp 1681620392
transform 1 0 2932 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4639
timestamp 1681620392
transform 1 0 2940 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4721
timestamp 1681620392
transform 1 0 2908 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4722
timestamp 1681620392
transform 1 0 2924 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4723
timestamp 1681620392
transform 1 0 2940 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_4062
timestamp 1681620392
transform 1 0 2924 0 1 595
box -3 -3 3 3
use Project_Top_VIA0  Project_Top_VIA0_48
timestamp 1681620392
transform 1 0 48 0 1 570
box -10 -3 10 3
use FILL  FILL_1180
timestamp 1681620392
transform 1 0 72 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_4079
timestamp 1681620392
transform 1 0 92 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_257
timestamp 1681620392
transform 1 0 80 0 1 570
box -8 -3 104 105
use INVX2  INVX2_304
timestamp 1681620392
transform 1 0 176 0 1 570
box -9 -3 26 105
use FILL  FILL_1182
timestamp 1681620392
transform 1 0 192 0 1 570
box -8 -3 16 105
use FILL  FILL_1191
timestamp 1681620392
transform 1 0 200 0 1 570
box -8 -3 16 105
use FILL  FILL_1193
timestamp 1681620392
transform 1 0 208 0 1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_90
timestamp 1681620392
transform 1 0 216 0 1 570
box -8 -3 32 105
use INVX2  INVX2_306
timestamp 1681620392
transform 1 0 240 0 1 570
box -9 -3 26 105
use FILL  FILL_1195
timestamp 1681620392
transform 1 0 256 0 1 570
box -8 -3 16 105
use FILL  FILL_1196
timestamp 1681620392
transform 1 0 264 0 1 570
box -8 -3 16 105
use FILL  FILL_1197
timestamp 1681620392
transform 1 0 272 0 1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_91
timestamp 1681620392
transform -1 0 304 0 1 570
box -8 -3 32 105
use FILL  FILL_1201
timestamp 1681620392
transform 1 0 304 0 1 570
box -8 -3 16 105
use FILL  FILL_1202
timestamp 1681620392
transform 1 0 312 0 1 570
box -8 -3 16 105
use AOI21X1  AOI21X1_32
timestamp 1681620392
transform 1 0 320 0 1 570
box -7 -3 39 105
use M3_M2  M3_M2_4080
timestamp 1681620392
transform 1 0 364 0 1 575
box -3 -3 3 3
use FILL  FILL_1203
timestamp 1681620392
transform 1 0 352 0 1 570
box -8 -3 16 105
use INVX2  INVX2_307
timestamp 1681620392
transform -1 0 376 0 1 570
box -9 -3 26 105
use NAND2X1  NAND2X1_268
timestamp 1681620392
transform -1 0 400 0 1 570
box -8 -3 32 105
use M3_M2  M3_M2_4081
timestamp 1681620392
transform 1 0 420 0 1 575
box -3 -3 3 3
use NAND2X1  NAND2X1_269
timestamp 1681620392
transform -1 0 424 0 1 570
box -8 -3 32 105
use NAND3X1  NAND3X1_97
timestamp 1681620392
transform 1 0 424 0 1 570
box -8 -3 40 105
use M3_M2  M3_M2_4082
timestamp 1681620392
transform 1 0 468 0 1 575
box -3 -3 3 3
use INVX2  INVX2_308
timestamp 1681620392
transform 1 0 456 0 1 570
box -9 -3 26 105
use NAND2X1  NAND2X1_270
timestamp 1681620392
transform -1 0 496 0 1 570
box -8 -3 32 105
use AOI21X1  AOI21X1_33
timestamp 1681620392
transform 1 0 496 0 1 570
box -7 -3 39 105
use FILL  FILL_1213
timestamp 1681620392
transform 1 0 528 0 1 570
box -8 -3 16 105
use FILL  FILL_1214
timestamp 1681620392
transform 1 0 536 0 1 570
box -8 -3 16 105
use FILL  FILL_1215
timestamp 1681620392
transform 1 0 544 0 1 570
box -8 -3 16 105
use INVX2  INVX2_309
timestamp 1681620392
transform 1 0 552 0 1 570
box -9 -3 26 105
use M3_M2  M3_M2_4083
timestamp 1681620392
transform 1 0 588 0 1 575
box -3 -3 3 3
use NAND2X1  NAND2X1_275
timestamp 1681620392
transform -1 0 592 0 1 570
box -8 -3 32 105
use FILL  FILL_1216
timestamp 1681620392
transform 1 0 592 0 1 570
box -8 -3 16 105
use FILL  FILL_1217
timestamp 1681620392
transform 1 0 600 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_4084
timestamp 1681620392
transform 1 0 644 0 1 575
box -3 -3 3 3
use OAI21X1  OAI21X1_268
timestamp 1681620392
transform 1 0 608 0 1 570
box -8 -3 34 105
use NAND2X1  NAND2X1_276
timestamp 1681620392
transform 1 0 640 0 1 570
box -8 -3 32 105
use OAI21X1  OAI21X1_269
timestamp 1681620392
transform 1 0 664 0 1 570
box -8 -3 34 105
use INVX2  INVX2_310
timestamp 1681620392
transform 1 0 696 0 1 570
box -9 -3 26 105
use OAI22X1  OAI22X1_95
timestamp 1681620392
transform -1 0 752 0 1 570
box -8 -3 46 105
use FILL  FILL_1220
timestamp 1681620392
transform 1 0 752 0 1 570
box -8 -3 16 105
use FILL  FILL_1221
timestamp 1681620392
transform 1 0 760 0 1 570
box -8 -3 16 105
use FILL  FILL_1222
timestamp 1681620392
transform 1 0 768 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_258
timestamp 1681620392
transform 1 0 776 0 1 570
box -8 -3 104 105
use INVX2  INVX2_311
timestamp 1681620392
transform -1 0 888 0 1 570
box -9 -3 26 105
use FILL  FILL_1223
timestamp 1681620392
transform 1 0 888 0 1 570
box -8 -3 16 105
use FILL  FILL_1224
timestamp 1681620392
transform 1 0 896 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_271
timestamp 1681620392
transform -1 0 936 0 1 570
box -8 -3 34 105
use M3_M2  M3_M2_4085
timestamp 1681620392
transform 1 0 988 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_259
timestamp 1681620392
transform 1 0 936 0 1 570
box -8 -3 104 105
use INVX2  INVX2_312
timestamp 1681620392
transform -1 0 1048 0 1 570
box -9 -3 26 105
use M3_M2  M3_M2_4086
timestamp 1681620392
transform 1 0 1084 0 1 575
box -3 -3 3 3
use OAI22X1  OAI22X1_96
timestamp 1681620392
transform 1 0 1048 0 1 570
box -8 -3 46 105
use FILL  FILL_1225
timestamp 1681620392
transform 1 0 1088 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_99
timestamp 1681620392
transform 1 0 1096 0 1 570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_262
timestamp 1681620392
transform -1 0 1232 0 1 570
box -8 -3 104 105
use BUFX2  BUFX2_38
timestamp 1681620392
transform -1 0 1256 0 1 570
box -5 -3 28 105
use FILL  FILL_1235
timestamp 1681620392
transform 1 0 1256 0 1 570
box -8 -3 16 105
use BUFX2  BUFX2_39
timestamp 1681620392
transform 1 0 1264 0 1 570
box -5 -3 28 105
use AOI21X1  AOI21X1_34
timestamp 1681620392
transform -1 0 1320 0 1 570
box -7 -3 39 105
use M3_M2  M3_M2_4087
timestamp 1681620392
transform 1 0 1348 0 1 575
box -3 -3 3 3
use NAND2X1  NAND2X1_279
timestamp 1681620392
transform 1 0 1320 0 1 570
box -8 -3 32 105
use INVX2  INVX2_315
timestamp 1681620392
transform 1 0 1344 0 1 570
box -9 -3 26 105
use AOI21X1  AOI21X1_35
timestamp 1681620392
transform 1 0 1360 0 1 570
box -7 -3 39 105
use OAI22X1  OAI22X1_100
timestamp 1681620392
transform 1 0 1392 0 1 570
box -8 -3 46 105
use AOI21X1  AOI21X1_36
timestamp 1681620392
transform -1 0 1464 0 1 570
box -7 -3 39 105
use OAI21X1  OAI21X1_272
timestamp 1681620392
transform -1 0 1496 0 1 570
box -8 -3 34 105
use INVX2  INVX2_316
timestamp 1681620392
transform -1 0 1512 0 1 570
box -9 -3 26 105
use AOI21X1  AOI21X1_37
timestamp 1681620392
transform -1 0 1544 0 1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_38
timestamp 1681620392
transform 1 0 1544 0 1 570
box -7 -3 39 105
use OAI21X1  OAI21X1_273
timestamp 1681620392
transform 1 0 1576 0 1 570
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_263
timestamp 1681620392
transform 1 0 1608 0 1 570
box -8 -3 104 105
use FILL  FILL_1236
timestamp 1681620392
transform 1 0 1704 0 1 570
box -8 -3 16 105
use INVX2  INVX2_317
timestamp 1681620392
transform -1 0 1728 0 1 570
box -9 -3 26 105
use FILL  FILL_1237
timestamp 1681620392
transform 1 0 1728 0 1 570
box -8 -3 16 105
use FILL  FILL_1238
timestamp 1681620392
transform 1 0 1736 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_101
timestamp 1681620392
transform -1 0 1784 0 1 570
box -8 -3 46 105
use M3_M2  M3_M2_4088
timestamp 1681620392
transform 1 0 1796 0 1 575
box -3 -3 3 3
use FILL  FILL_1239
timestamp 1681620392
transform 1 0 1784 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_264
timestamp 1681620392
transform 1 0 1792 0 1 570
box -8 -3 104 105
use FILL  FILL_1240
timestamp 1681620392
transform 1 0 1888 0 1 570
box -8 -3 16 105
use INVX2  INVX2_318
timestamp 1681620392
transform 1 0 1896 0 1 570
box -9 -3 26 105
use OAI21X1  OAI21X1_274
timestamp 1681620392
transform 1 0 1912 0 1 570
box -8 -3 34 105
use NAND2X1  NAND2X1_280
timestamp 1681620392
transform -1 0 1968 0 1 570
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_265
timestamp 1681620392
transform 1 0 1968 0 1 570
box -8 -3 104 105
use NAND2X1  NAND2X1_281
timestamp 1681620392
transform 1 0 2064 0 1 570
box -8 -3 32 105
use M3_M2  M3_M2_4089
timestamp 1681620392
transform 1 0 2132 0 1 575
box -3 -3 3 3
use OAI22X1  OAI22X1_102
timestamp 1681620392
transform -1 0 2128 0 1 570
box -8 -3 46 105
use M3_M2  M3_M2_4090
timestamp 1681620392
transform 1 0 2188 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_266
timestamp 1681620392
transform 1 0 2128 0 1 570
box -8 -3 104 105
use INVX2  INVX2_319
timestamp 1681620392
transform 1 0 2224 0 1 570
box -9 -3 26 105
use M3_M2  M3_M2_4091
timestamp 1681620392
transform 1 0 2276 0 1 575
box -3 -3 3 3
use OAI21X1  OAI21X1_275
timestamp 1681620392
transform 1 0 2240 0 1 570
box -8 -3 34 105
use NAND2X1  NAND2X1_282
timestamp 1681620392
transform -1 0 2296 0 1 570
box -8 -3 32 105
use M3_M2  M3_M2_4092
timestamp 1681620392
transform 1 0 2316 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_267
timestamp 1681620392
transform 1 0 2296 0 1 570
box -8 -3 104 105
use NAND2X1  NAND2X1_283
timestamp 1681620392
transform 1 0 2392 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_284
timestamp 1681620392
transform 1 0 2416 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_285
timestamp 1681620392
transform 1 0 2440 0 1 570
box -8 -3 32 105
use FILL  FILL_1241
timestamp 1681620392
transform 1 0 2464 0 1 570
box -8 -3 16 105
use FILL  FILL_1242
timestamp 1681620392
transform 1 0 2472 0 1 570
box -8 -3 16 105
use FILL  FILL_1243
timestamp 1681620392
transform 1 0 2480 0 1 570
box -8 -3 16 105
use INVX2  INVX2_320
timestamp 1681620392
transform -1 0 2504 0 1 570
box -9 -3 26 105
use FILL  FILL_1244
timestamp 1681620392
transform 1 0 2504 0 1 570
box -8 -3 16 105
use FILL  FILL_1245
timestamp 1681620392
transform 1 0 2512 0 1 570
box -8 -3 16 105
use FILL  FILL_1246
timestamp 1681620392
transform 1 0 2520 0 1 570
box -8 -3 16 105
use FILL  FILL_1247
timestamp 1681620392
transform 1 0 2528 0 1 570
box -8 -3 16 105
use FILL  FILL_1248
timestamp 1681620392
transform 1 0 2536 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_276
timestamp 1681620392
transform -1 0 2576 0 1 570
box -8 -3 34 105
use FILL  FILL_1249
timestamp 1681620392
transform 1 0 2576 0 1 570
box -8 -3 16 105
use FILL  FILL_1250
timestamp 1681620392
transform 1 0 2584 0 1 570
box -8 -3 16 105
use FILL  FILL_1251
timestamp 1681620392
transform 1 0 2592 0 1 570
box -8 -3 16 105
use FILL  FILL_1252
timestamp 1681620392
transform 1 0 2600 0 1 570
box -8 -3 16 105
use FILL  FILL_1253
timestamp 1681620392
transform 1 0 2608 0 1 570
box -8 -3 16 105
use INVX2  INVX2_321
timestamp 1681620392
transform -1 0 2632 0 1 570
box -9 -3 26 105
use FILL  FILL_1254
timestamp 1681620392
transform 1 0 2632 0 1 570
box -8 -3 16 105
use FILL  FILL_1255
timestamp 1681620392
transform 1 0 2640 0 1 570
box -8 -3 16 105
use FILL  FILL_1256
timestamp 1681620392
transform 1 0 2648 0 1 570
box -8 -3 16 105
use FILL  FILL_1257
timestamp 1681620392
transform 1 0 2656 0 1 570
box -8 -3 16 105
use FILL  FILL_1258
timestamp 1681620392
transform 1 0 2664 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_277
timestamp 1681620392
transform -1 0 2704 0 1 570
box -8 -3 34 105
use FILL  FILL_1259
timestamp 1681620392
transform 1 0 2704 0 1 570
box -8 -3 16 105
use INVX2  INVX2_322
timestamp 1681620392
transform -1 0 2728 0 1 570
box -9 -3 26 105
use FILL  FILL_1260
timestamp 1681620392
transform 1 0 2728 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_268
timestamp 1681620392
transform -1 0 2832 0 1 570
box -8 -3 104 105
use FILL  FILL_1261
timestamp 1681620392
transform 1 0 2832 0 1 570
box -8 -3 16 105
use FILL  FILL_1262
timestamp 1681620392
transform 1 0 2840 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_43
timestamp 1681620392
transform -1 0 2888 0 1 570
box -8 -3 46 105
use FILL  FILL_1263
timestamp 1681620392
transform 1 0 2888 0 1 570
box -8 -3 16 105
use FILL  FILL_1264
timestamp 1681620392
transform 1 0 2896 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_103
timestamp 1681620392
transform -1 0 2944 0 1 570
box -8 -3 46 105
use FILL  FILL_1265
timestamp 1681620392
transform 1 0 2944 0 1 570
box -8 -3 16 105
use FILL  FILL_1266
timestamp 1681620392
transform 1 0 2952 0 1 570
box -8 -3 16 105
use FILL  FILL_1267
timestamp 1681620392
transform 1 0 2960 0 1 570
box -8 -3 16 105
use FILL  FILL_1300
timestamp 1681620392
transform 1 0 2968 0 1 570
box -8 -3 16 105
use FILL  FILL_1302
timestamp 1681620392
transform 1 0 2976 0 1 570
box -8 -3 16 105
use INVX2  INVX2_332
timestamp 1681620392
transform 1 0 2984 0 1 570
box -9 -3 26 105
use FILL  FILL_1304
timestamp 1681620392
transform 1 0 3000 0 1 570
box -8 -3 16 105
use FILL  FILL_1308
timestamp 1681620392
transform 1 0 3008 0 1 570
box -8 -3 16 105
use Project_Top_VIA0  Project_Top_VIA0_49
timestamp 1681620392
transform 1 0 3043 0 1 570
box -10 -3 10 3
use M3_M2  M3_M2_4200
timestamp 1681620392
transform 1 0 116 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_4735
timestamp 1681620392
transform 1 0 124 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_4128
timestamp 1681620392
transform 1 0 164 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4156
timestamp 1681620392
transform 1 0 140 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_4736
timestamp 1681620392
transform 1 0 148 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_4157
timestamp 1681620392
transform 1 0 156 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_4737
timestamp 1681620392
transform 1 0 164 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4738
timestamp 1681620392
transform 1 0 172 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4818
timestamp 1681620392
transform 1 0 140 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4819
timestamp 1681620392
transform 1 0 156 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4820
timestamp 1681620392
transform 1 0 164 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4201
timestamp 1681620392
transform 1 0 156 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4202
timestamp 1681620392
transform 1 0 172 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4129
timestamp 1681620392
transform 1 0 188 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4105
timestamp 1681620392
transform 1 0 268 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_4739
timestamp 1681620392
transform 1 0 252 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4740
timestamp 1681620392
transform 1 0 268 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4821
timestamp 1681620392
transform 1 0 244 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4822
timestamp 1681620392
transform 1 0 260 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4203
timestamp 1681620392
transform 1 0 260 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_4823
timestamp 1681620392
transform 1 0 276 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4106
timestamp 1681620392
transform 1 0 300 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_4733
timestamp 1681620392
transform 1 0 300 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_4130
timestamp 1681620392
transform 1 0 308 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4741
timestamp 1681620392
transform 1 0 308 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4742
timestamp 1681620392
transform 1 0 316 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4743
timestamp 1681620392
transform 1 0 332 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4824
timestamp 1681620392
transform 1 0 324 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4228
timestamp 1681620392
transform 1 0 316 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4131
timestamp 1681620392
transform 1 0 372 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4744
timestamp 1681620392
transform 1 0 388 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4825
timestamp 1681620392
transform 1 0 396 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4177
timestamp 1681620392
transform 1 0 404 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_4894
timestamp 1681620392
transform 1 0 388 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_4229
timestamp 1681620392
transform 1 0 388 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_4826
timestamp 1681620392
transform 1 0 420 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4895
timestamp 1681620392
transform 1 0 412 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_4204
timestamp 1681620392
transform 1 0 420 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4132
timestamp 1681620392
transform 1 0 444 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4158
timestamp 1681620392
transform 1 0 436 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_4745
timestamp 1681620392
transform 1 0 444 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4827
timestamp 1681620392
transform 1 0 436 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4746
timestamp 1681620392
transform 1 0 468 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4747
timestamp 1681620392
transform 1 0 484 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4828
timestamp 1681620392
transform 1 0 492 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4896
timestamp 1681620392
transform 1 0 484 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_4230
timestamp 1681620392
transform 1 0 492 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_4829
timestamp 1681620392
transform 1 0 508 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4178
timestamp 1681620392
transform 1 0 516 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_4830
timestamp 1681620392
transform 1 0 524 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4179
timestamp 1681620392
transform 1 0 532 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_4748
timestamp 1681620392
transform 1 0 564 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4831
timestamp 1681620392
transform 1 0 540 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4205
timestamp 1681620392
transform 1 0 508 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4180
timestamp 1681620392
transform 1 0 564 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_4897
timestamp 1681620392
transform 1 0 540 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4898
timestamp 1681620392
transform 1 0 564 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4919
timestamp 1681620392
transform 1 0 532 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_4749
timestamp 1681620392
transform 1 0 580 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_4159
timestamp 1681620392
transform 1 0 588 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4181
timestamp 1681620392
transform 1 0 580 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4093
timestamp 1681620392
transform 1 0 620 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_4750
timestamp 1681620392
transform 1 0 620 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4751
timestamp 1681620392
transform 1 0 628 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4832
timestamp 1681620392
transform 1 0 596 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4833
timestamp 1681620392
transform 1 0 604 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4899
timestamp 1681620392
transform 1 0 588 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_4231
timestamp 1681620392
transform 1 0 580 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4243
timestamp 1681620392
transform 1 0 572 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4244
timestamp 1681620392
transform 1 0 596 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4160
timestamp 1681620392
transform 1 0 660 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_4834
timestamp 1681620392
transform 1 0 636 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4835
timestamp 1681620392
transform 1 0 652 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4900
timestamp 1681620392
transform 1 0 628 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_4206
timestamp 1681620392
transform 1 0 636 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_4901
timestamp 1681620392
transform 1 0 660 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4920
timestamp 1681620392
transform 1 0 668 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_4921
timestamp 1681620392
transform 1 0 684 0 1 505
box -2 -2 2 2
use M3_M2  M3_M2_4107
timestamp 1681620392
transform 1 0 708 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4133
timestamp 1681620392
transform 1 0 700 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4902
timestamp 1681620392
transform 1 0 700 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_4245
timestamp 1681620392
transform 1 0 692 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_4903
timestamp 1681620392
transform 1 0 724 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_4246
timestamp 1681620392
transform 1 0 724 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4108
timestamp 1681620392
transform 1 0 748 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4134
timestamp 1681620392
transform 1 0 756 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4135
timestamp 1681620392
transform 1 0 772 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4752
timestamp 1681620392
transform 1 0 748 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4753
timestamp 1681620392
transform 1 0 756 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4754
timestamp 1681620392
transform 1 0 772 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4755
timestamp 1681620392
transform 1 0 788 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4836
timestamp 1681620392
transform 1 0 748 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4837
timestamp 1681620392
transform 1 0 764 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4207
timestamp 1681620392
transform 1 0 788 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4232
timestamp 1681620392
transform 1 0 796 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_4756
timestamp 1681620392
transform 1 0 820 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_4161
timestamp 1681620392
transform 1 0 828 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_4838
timestamp 1681620392
transform 1 0 820 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4208
timestamp 1681620392
transform 1 0 820 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4094
timestamp 1681620392
transform 1 0 852 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4136
timestamp 1681620392
transform 1 0 876 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4095
timestamp 1681620392
transform 1 0 948 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4137
timestamp 1681620392
transform 1 0 948 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4138
timestamp 1681620392
transform 1 0 980 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4757
timestamp 1681620392
transform 1 0 836 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4758
timestamp 1681620392
transform 1 0 852 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_4162
timestamp 1681620392
transform 1 0 932 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4096
timestamp 1681620392
transform 1 0 1052 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_4759
timestamp 1681620392
transform 1 0 948 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_4182
timestamp 1681620392
transform 1 0 836 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_4839
timestamp 1681620392
transform 1 0 876 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4183
timestamp 1681620392
transform 1 0 884 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4163
timestamp 1681620392
transform 1 0 1028 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_4760
timestamp 1681620392
transform 1 0 1036 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_4164
timestamp 1681620392
transform 1 0 1044 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4109
timestamp 1681620392
transform 1 0 1084 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4139
timestamp 1681620392
transform 1 0 1076 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4761
timestamp 1681620392
transform 1 0 1052 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4762
timestamp 1681620392
transform 1 0 1068 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4840
timestamp 1681620392
transform 1 0 932 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4841
timestamp 1681620392
transform 1 0 972 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4233
timestamp 1681620392
transform 1 0 844 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4184
timestamp 1681620392
transform 1 0 1020 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_4842
timestamp 1681620392
transform 1 0 1028 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4843
timestamp 1681620392
transform 1 0 1036 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4844
timestamp 1681620392
transform 1 0 1044 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4845
timestamp 1681620392
transform 1 0 1060 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4185
timestamp 1681620392
transform 1 0 1068 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4209
timestamp 1681620392
transform 1 0 1012 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4210
timestamp 1681620392
transform 1 0 1028 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4211
timestamp 1681620392
transform 1 0 1044 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4247
timestamp 1681620392
transform 1 0 948 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4234
timestamp 1681620392
transform 1 0 1060 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_4904
timestamp 1681620392
transform 1 0 1084 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_4110
timestamp 1681620392
transform 1 0 1124 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_4763
timestamp 1681620392
transform 1 0 1108 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_4140
timestamp 1681620392
transform 1 0 1132 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4764
timestamp 1681620392
transform 1 0 1132 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4765
timestamp 1681620392
transform 1 0 1156 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_4165
timestamp 1681620392
transform 1 0 1164 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_4766
timestamp 1681620392
transform 1 0 1180 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4767
timestamp 1681620392
transform 1 0 1196 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4846
timestamp 1681620392
transform 1 0 1164 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4847
timestamp 1681620392
transform 1 0 1188 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4848
timestamp 1681620392
transform 1 0 1204 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4235
timestamp 1681620392
transform 1 0 1188 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4111
timestamp 1681620392
transform 1 0 1324 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4141
timestamp 1681620392
transform 1 0 1284 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4768
timestamp 1681620392
transform 1 0 1220 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4769
timestamp 1681620392
transform 1 0 1236 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_4258
timestamp 1681620392
transform 1 0 1204 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4166
timestamp 1681620392
transform 1 0 1308 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_4770
timestamp 1681620392
transform 1 0 1324 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_4167
timestamp 1681620392
transform 1 0 1332 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_4771
timestamp 1681620392
transform 1 0 1348 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4849
timestamp 1681620392
transform 1 0 1284 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4850
timestamp 1681620392
transform 1 0 1316 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4851
timestamp 1681620392
transform 1 0 1332 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4852
timestamp 1681620392
transform 1 0 1348 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4212
timestamp 1681620392
transform 1 0 1300 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4248
timestamp 1681620392
transform 1 0 1236 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4249
timestamp 1681620392
transform 1 0 1260 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4259
timestamp 1681620392
transform 1 0 1284 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4186
timestamp 1681620392
transform 1 0 1356 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4213
timestamp 1681620392
transform 1 0 1332 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_4905
timestamp 1681620392
transform 1 0 1348 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4772
timestamp 1681620392
transform 1 0 1372 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4906
timestamp 1681620392
transform 1 0 1372 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_4097
timestamp 1681620392
transform 1 0 1388 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4168
timestamp 1681620392
transform 1 0 1396 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_4853
timestamp 1681620392
transform 1 0 1396 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4214
timestamp 1681620392
transform 1 0 1396 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_4922
timestamp 1681620392
transform 1 0 1396 0 1 505
box -2 -2 2 2
use M3_M2  M3_M2_4142
timestamp 1681620392
transform 1 0 1412 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4143
timestamp 1681620392
transform 1 0 1428 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4773
timestamp 1681620392
transform 1 0 1428 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4854
timestamp 1681620392
transform 1 0 1420 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4187
timestamp 1681620392
transform 1 0 1428 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4098
timestamp 1681620392
transform 1 0 1468 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4099
timestamp 1681620392
transform 1 0 1500 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4112
timestamp 1681620392
transform 1 0 1492 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4144
timestamp 1681620392
transform 1 0 1484 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4774
timestamp 1681620392
transform 1 0 1476 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4855
timestamp 1681620392
transform 1 0 1452 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4856
timestamp 1681620392
transform 1 0 1460 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4215
timestamp 1681620392
transform 1 0 1436 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4188
timestamp 1681620392
transform 1 0 1468 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_4857
timestamp 1681620392
transform 1 0 1476 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4907
timestamp 1681620392
transform 1 0 1444 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_4236
timestamp 1681620392
transform 1 0 1444 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_4908
timestamp 1681620392
transform 1 0 1476 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_4169
timestamp 1681620392
transform 1 0 1492 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_4909
timestamp 1681620392
transform 1 0 1492 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4858
timestamp 1681620392
transform 1 0 1524 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4775
timestamp 1681620392
transform 1 0 1548 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4859
timestamp 1681620392
transform 1 0 1556 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4145
timestamp 1681620392
transform 1 0 1564 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4776
timestamp 1681620392
transform 1 0 1564 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4860
timestamp 1681620392
transform 1 0 1564 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4216
timestamp 1681620392
transform 1 0 1556 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4237
timestamp 1681620392
transform 1 0 1564 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4113
timestamp 1681620392
transform 1 0 1580 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4114
timestamp 1681620392
transform 1 0 1604 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_4777
timestamp 1681620392
transform 1 0 1580 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4778
timestamp 1681620392
transform 1 0 1588 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4861
timestamp 1681620392
transform 1 0 1580 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4217
timestamp 1681620392
transform 1 0 1580 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4115
timestamp 1681620392
transform 1 0 1620 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4238
timestamp 1681620392
transform 1 0 1612 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_4910
timestamp 1681620392
transform 1 0 1620 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4779
timestamp 1681620392
transform 1 0 1636 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_4218
timestamp 1681620392
transform 1 0 1636 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4116
timestamp 1681620392
transform 1 0 1652 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4146
timestamp 1681620392
transform 1 0 1732 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4780
timestamp 1681620392
transform 1 0 1652 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4862
timestamp 1681620392
transform 1 0 1676 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4189
timestamp 1681620392
transform 1 0 1692 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_4781
timestamp 1681620392
transform 1 0 1740 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4863
timestamp 1681620392
transform 1 0 1732 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4219
timestamp 1681620392
transform 1 0 1676 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4190
timestamp 1681620392
transform 1 0 1740 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4117
timestamp 1681620392
transform 1 0 1780 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_4782
timestamp 1681620392
transform 1 0 1772 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4783
timestamp 1681620392
transform 1 0 1788 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4784
timestamp 1681620392
transform 1 0 1804 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4864
timestamp 1681620392
transform 1 0 1780 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4865
timestamp 1681620392
transform 1 0 1796 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4866
timestamp 1681620392
transform 1 0 1812 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4250
timestamp 1681620392
transform 1 0 1804 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_4785
timestamp 1681620392
transform 1 0 1836 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4786
timestamp 1681620392
transform 1 0 1844 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4787
timestamp 1681620392
transform 1 0 1884 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4867
timestamp 1681620392
transform 1 0 1860 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4220
timestamp 1681620392
transform 1 0 1860 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4118
timestamp 1681620392
transform 1 0 1924 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4100
timestamp 1681620392
transform 1 0 1964 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4101
timestamp 1681620392
transform 1 0 2036 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4147
timestamp 1681620392
transform 1 0 1940 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4148
timestamp 1681620392
transform 1 0 1980 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4788
timestamp 1681620392
transform 1 0 1908 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4789
timestamp 1681620392
transform 1 0 1916 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4790
timestamp 1681620392
transform 1 0 1940 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4791
timestamp 1681620392
transform 1 0 1956 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4792
timestamp 1681620392
transform 1 0 2044 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4793
timestamp 1681620392
transform 1 0 2060 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4794
timestamp 1681620392
transform 1 0 2076 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4795
timestamp 1681620392
transform 1 0 2084 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4868
timestamp 1681620392
transform 1 0 1892 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4191
timestamp 1681620392
transform 1 0 1908 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_4869
timestamp 1681620392
transform 1 0 1924 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4221
timestamp 1681620392
transform 1 0 1892 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4251
timestamp 1681620392
transform 1 0 1876 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_4870
timestamp 1681620392
transform 1 0 1980 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4871
timestamp 1681620392
transform 1 0 2036 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4872
timestamp 1681620392
transform 1 0 2052 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4911
timestamp 1681620392
transform 1 0 1940 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_4252
timestamp 1681620392
transform 1 0 1900 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4253
timestamp 1681620392
transform 1 0 1916 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4149
timestamp 1681620392
transform 1 0 2116 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4796
timestamp 1681620392
transform 1 0 2100 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_4170
timestamp 1681620392
transform 1 0 2108 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4119
timestamp 1681620392
transform 1 0 2148 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4150
timestamp 1681620392
transform 1 0 2172 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4797
timestamp 1681620392
transform 1 0 2116 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4798
timestamp 1681620392
transform 1 0 2132 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4799
timestamp 1681620392
transform 1 0 2148 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_4171
timestamp 1681620392
transform 1 0 2180 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_4873
timestamp 1681620392
transform 1 0 2092 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4874
timestamp 1681620392
transform 1 0 2108 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4875
timestamp 1681620392
transform 1 0 2132 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4192
timestamp 1681620392
transform 1 0 2148 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_4876
timestamp 1681620392
transform 1 0 2172 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4222
timestamp 1681620392
transform 1 0 2132 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4260
timestamp 1681620392
transform 1 0 2204 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4120
timestamp 1681620392
transform 1 0 2268 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_4800
timestamp 1681620392
transform 1 0 2252 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4877
timestamp 1681620392
transform 1 0 2244 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4223
timestamp 1681620392
transform 1 0 2244 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4261
timestamp 1681620392
transform 1 0 2252 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4102
timestamp 1681620392
transform 1 0 2380 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4121
timestamp 1681620392
transform 1 0 2292 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4122
timestamp 1681620392
transform 1 0 2308 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4123
timestamp 1681620392
transform 1 0 2332 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_4801
timestamp 1681620392
transform 1 0 2276 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4802
timestamp 1681620392
transform 1 0 2292 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4803
timestamp 1681620392
transform 1 0 2380 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_4193
timestamp 1681620392
transform 1 0 2276 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_4878
timestamp 1681620392
transform 1 0 2316 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4194
timestamp 1681620392
transform 1 0 2356 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_4879
timestamp 1681620392
transform 1 0 2372 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4912
timestamp 1681620392
transform 1 0 2276 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4804
timestamp 1681620392
transform 1 0 2396 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_4103
timestamp 1681620392
transform 1 0 2452 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4124
timestamp 1681620392
transform 1 0 2444 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4151
timestamp 1681620392
transform 1 0 2428 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4805
timestamp 1681620392
transform 1 0 2428 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4880
timestamp 1681620392
transform 1 0 2404 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4881
timestamp 1681620392
transform 1 0 2420 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4125
timestamp 1681620392
transform 1 0 2492 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4152
timestamp 1681620392
transform 1 0 2492 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4806
timestamp 1681620392
transform 1 0 2452 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4807
timestamp 1681620392
transform 1 0 2468 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4882
timestamp 1681620392
transform 1 0 2444 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4913
timestamp 1681620392
transform 1 0 2396 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4914
timestamp 1681620392
transform 1 0 2420 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4915
timestamp 1681620392
transform 1 0 2428 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_4239
timestamp 1681620392
transform 1 0 2404 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4240
timestamp 1681620392
transform 1 0 2428 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4254
timestamp 1681620392
transform 1 0 2412 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4255
timestamp 1681620392
transform 1 0 2444 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4195
timestamp 1681620392
transform 1 0 2468 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4104
timestamp 1681620392
transform 1 0 2564 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4172
timestamp 1681620392
transform 1 0 2556 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_4883
timestamp 1681620392
transform 1 0 2492 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4884
timestamp 1681620392
transform 1 0 2548 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4256
timestamp 1681620392
transform 1 0 2564 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_4808
timestamp 1681620392
transform 1 0 2580 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_4173
timestamp 1681620392
transform 1 0 2604 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4174
timestamp 1681620392
transform 1 0 2652 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4196
timestamp 1681620392
transform 1 0 2580 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_4885
timestamp 1681620392
transform 1 0 2604 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4197
timestamp 1681620392
transform 1 0 2628 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_4886
timestamp 1681620392
transform 1 0 2660 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4224
timestamp 1681620392
transform 1 0 2620 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4257
timestamp 1681620392
transform 1 0 2596 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4175
timestamp 1681620392
transform 1 0 2684 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_4809
timestamp 1681620392
transform 1 0 2708 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4887
timestamp 1681620392
transform 1 0 2684 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4888
timestamp 1681620392
transform 1 0 2700 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4198
timestamp 1681620392
transform 1 0 2708 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4225
timestamp 1681620392
transform 1 0 2684 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4226
timestamp 1681620392
transform 1 0 2700 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_4889
timestamp 1681620392
transform 1 0 2724 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4916
timestamp 1681620392
transform 1 0 2724 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_4176
timestamp 1681620392
transform 1 0 2740 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_4917
timestamp 1681620392
transform 1 0 2740 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4890
timestamp 1681620392
transform 1 0 2756 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4153
timestamp 1681620392
transform 1 0 2780 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4810
timestamp 1681620392
transform 1 0 2780 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4811
timestamp 1681620392
transform 1 0 2788 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_4227
timestamp 1681620392
transform 1 0 2788 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_4812
timestamp 1681620392
transform 1 0 2844 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4734
timestamp 1681620392
transform 1 0 2860 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_4126
timestamp 1681620392
transform 1 0 2876 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_4813
timestamp 1681620392
transform 1 0 2876 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4814
timestamp 1681620392
transform 1 0 2884 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4891
timestamp 1681620392
transform 1 0 2892 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4918
timestamp 1681620392
transform 1 0 2908 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_4127
timestamp 1681620392
transform 1 0 2940 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4154
timestamp 1681620392
transform 1 0 2932 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4155
timestamp 1681620392
transform 1 0 2948 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_4815
timestamp 1681620392
transform 1 0 2916 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4816
timestamp 1681620392
transform 1 0 2940 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4817
timestamp 1681620392
transform 1 0 2956 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4892
timestamp 1681620392
transform 1 0 2932 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4893
timestamp 1681620392
transform 1 0 2940 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_4241
timestamp 1681620392
transform 1 0 2908 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4199
timestamp 1681620392
transform 1 0 2948 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4242
timestamp 1681620392
transform 1 0 2940 0 1 505
box -3 -3 3 3
use Project_Top_VIA0  Project_Top_VIA0_50
timestamp 1681620392
transform 1 0 24 0 1 470
box -10 -3 10 3
use FILL  FILL_1181
timestamp 1681620392
transform 1 0 72 0 -1 570
box -8 -3 16 105
use FILL  FILL_1183
timestamp 1681620392
transform 1 0 80 0 -1 570
box -8 -3 16 105
use FILL  FILL_1184
timestamp 1681620392
transform 1 0 88 0 -1 570
box -8 -3 16 105
use FILL  FILL_1185
timestamp 1681620392
transform 1 0 96 0 -1 570
box -8 -3 16 105
use FILL  FILL_1186
timestamp 1681620392
transform 1 0 104 0 -1 570
box -8 -3 16 105
use FILL  FILL_1187
timestamp 1681620392
transform 1 0 112 0 -1 570
box -8 -3 16 105
use FILL  FILL_1188
timestamp 1681620392
transform 1 0 120 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_4262
timestamp 1681620392
transform 1 0 172 0 1 475
box -3 -3 3 3
use OAI22X1  OAI22X1_93
timestamp 1681620392
transform -1 0 168 0 -1 570
box -8 -3 46 105
use INVX2  INVX2_305
timestamp 1681620392
transform 1 0 168 0 -1 570
box -9 -3 26 105
use FILL  FILL_1189
timestamp 1681620392
transform 1 0 184 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_4263
timestamp 1681620392
transform 1 0 204 0 1 475
box -3 -3 3 3
use FILL  FILL_1190
timestamp 1681620392
transform 1 0 192 0 -1 570
box -8 -3 16 105
use FILL  FILL_1192
timestamp 1681620392
transform 1 0 200 0 -1 570
box -8 -3 16 105
use FILL  FILL_1194
timestamp 1681620392
transform 1 0 208 0 -1 570
box -8 -3 16 105
use FILL  FILL_1198
timestamp 1681620392
transform 1 0 216 0 -1 570
box -8 -3 16 105
use FILL  FILL_1199
timestamp 1681620392
transform 1 0 224 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_94
timestamp 1681620392
transform -1 0 272 0 -1 570
box -8 -3 46 105
use FILL  FILL_1200
timestamp 1681620392
transform 1 0 272 0 -1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_92
timestamp 1681620392
transform -1 0 304 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_93
timestamp 1681620392
transform 1 0 304 0 -1 570
box -8 -3 32 105
use FILL  FILL_1204
timestamp 1681620392
transform 1 0 328 0 -1 570
box -8 -3 16 105
use FILL  FILL_1205
timestamp 1681620392
transform 1 0 336 0 -1 570
box -8 -3 16 105
use FILL  FILL_1206
timestamp 1681620392
transform 1 0 344 0 -1 570
box -8 -3 16 105
use FILL  FILL_1207
timestamp 1681620392
transform 1 0 352 0 -1 570
box -8 -3 16 105
use FILL  FILL_1208
timestamp 1681620392
transform 1 0 360 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_271
timestamp 1681620392
transform 1 0 368 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_272
timestamp 1681620392
transform 1 0 392 0 -1 570
box -8 -3 32 105
use FILL  FILL_1209
timestamp 1681620392
transform 1 0 416 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_273
timestamp 1681620392
transform -1 0 448 0 -1 570
box -8 -3 32 105
use FILL  FILL_1210
timestamp 1681620392
transform 1 0 448 0 -1 570
box -8 -3 16 105
use FILL  FILL_1211
timestamp 1681620392
transform 1 0 456 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_274
timestamp 1681620392
transform 1 0 464 0 -1 570
box -8 -3 32 105
use FILL  FILL_1212
timestamp 1681620392
transform 1 0 488 0 -1 570
box -8 -3 16 105
use AND2X2  AND2X2_25
timestamp 1681620392
transform 1 0 496 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_98
timestamp 1681620392
transform 1 0 528 0 -1 570
box -8 -3 40 105
use NAND2X1  NAND2X1_277
timestamp 1681620392
transform 1 0 560 0 -1 570
box -8 -3 32 105
use FILL  FILL_1218
timestamp 1681620392
transform 1 0 584 0 -1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_270
timestamp 1681620392
transform 1 0 592 0 -1 570
box -8 -3 34 105
use AND2X2  AND2X2_26
timestamp 1681620392
transform 1 0 624 0 -1 570
box -8 -3 40 105
use FILL  FILL_1219
timestamp 1681620392
transform 1 0 656 0 -1 570
box -8 -3 16 105
use NAND3X1  NAND3X1_99
timestamp 1681620392
transform 1 0 664 0 -1 570
box -8 -3 40 105
use FILL  FILL_1226
timestamp 1681620392
transform 1 0 696 0 -1 570
box -8 -3 16 105
use FILL  FILL_1227
timestamp 1681620392
transform 1 0 704 0 -1 570
box -8 -3 16 105
use FILL  FILL_1228
timestamp 1681620392
transform 1 0 712 0 -1 570
box -8 -3 16 105
use FILL  FILL_1229
timestamp 1681620392
transform 1 0 720 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_278
timestamp 1681620392
transform -1 0 752 0 -1 570
box -8 -3 32 105
use OAI22X1  OAI22X1_97
timestamp 1681620392
transform -1 0 792 0 -1 570
box -8 -3 46 105
use FILL  FILL_1230
timestamp 1681620392
transform 1 0 792 0 -1 570
box -8 -3 16 105
use FILL  FILL_1231
timestamp 1681620392
transform 1 0 800 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_313
timestamp 1681620392
transform -1 0 824 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_314
timestamp 1681620392
transform -1 0 840 0 -1 570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_260
timestamp 1681620392
transform 1 0 840 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_261
timestamp 1681620392
transform 1 0 936 0 -1 570
box -8 -3 104 105
use OAI22X1  OAI22X1_98
timestamp 1681620392
transform 1 0 1032 0 -1 570
box -8 -3 46 105
use FILL  FILL_1232
timestamp 1681620392
transform 1 0 1072 0 -1 570
box -8 -3 16 105
use FILL  FILL_1233
timestamp 1681620392
transform 1 0 1080 0 -1 570
box -8 -3 16 105
use FILL  FILL_1234
timestamp 1681620392
transform 1 0 1088 0 -1 570
box -8 -3 16 105
use FILL  FILL_1268
timestamp 1681620392
transform 1 0 1096 0 -1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_278
timestamp 1681620392
transform -1 0 1136 0 -1 570
box -8 -3 34 105
use FILL  FILL_1269
timestamp 1681620392
transform 1 0 1136 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_323
timestamp 1681620392
transform -1 0 1160 0 -1 570
box -9 -3 26 105
use OAI22X1  OAI22X1_104
timestamp 1681620392
transform 1 0 1160 0 -1 570
box -8 -3 46 105
use BUFX2  BUFX2_40
timestamp 1681620392
transform 1 0 1200 0 -1 570
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_269
timestamp 1681620392
transform 1 0 1224 0 -1 570
box -8 -3 104 105
use OAI21X1  OAI21X1_279
timestamp 1681620392
transform 1 0 1320 0 -1 570
box -8 -3 34 105
use INVX2  INVX2_324
timestamp 1681620392
transform -1 0 1368 0 -1 570
box -9 -3 26 105
use FILL  FILL_1270
timestamp 1681620392
transform 1 0 1368 0 -1 570
box -8 -3 16 105
use NAND3X1  NAND3X1_100
timestamp 1681620392
transform -1 0 1408 0 -1 570
box -8 -3 40 105
use FILL  FILL_1271
timestamp 1681620392
transform 1 0 1408 0 -1 570
box -8 -3 16 105
use FILL  FILL_1272
timestamp 1681620392
transform 1 0 1416 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_286
timestamp 1681620392
transform 1 0 1424 0 -1 570
box -8 -3 32 105
use OAI21X1  OAI21X1_280
timestamp 1681620392
transform 1 0 1448 0 -1 570
box -8 -3 34 105
use FILL  FILL_1273
timestamp 1681620392
transform 1 0 1480 0 -1 570
box -8 -3 16 105
use FILL  FILL_1274
timestamp 1681620392
transform 1 0 1488 0 -1 570
box -8 -3 16 105
use FILL  FILL_1275
timestamp 1681620392
transform 1 0 1496 0 -1 570
box -8 -3 16 105
use AND2X2  AND2X2_27
timestamp 1681620392
transform -1 0 1536 0 -1 570
box -8 -3 40 105
use FILL  FILL_1276
timestamp 1681620392
transform 1 0 1536 0 -1 570
box -8 -3 16 105
use FILL  FILL_1277
timestamp 1681620392
transform 1 0 1544 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_325
timestamp 1681620392
transform -1 0 1568 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_326
timestamp 1681620392
transform -1 0 1584 0 -1 570
box -9 -3 26 105
use OAI21X1  OAI21X1_281
timestamp 1681620392
transform 1 0 1584 0 -1 570
box -8 -3 34 105
use FILL  FILL_1278
timestamp 1681620392
transform 1 0 1616 0 -1 570
box -8 -3 16 105
use FILL  FILL_1279
timestamp 1681620392
transform 1 0 1624 0 -1 570
box -8 -3 16 105
use FILL  FILL_1280
timestamp 1681620392
transform 1 0 1632 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_270
timestamp 1681620392
transform 1 0 1640 0 -1 570
box -8 -3 104 105
use FILL  FILL_1281
timestamp 1681620392
transform 1 0 1736 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_327
timestamp 1681620392
transform 1 0 1744 0 -1 570
box -9 -3 26 105
use FILL  FILL_1282
timestamp 1681620392
transform 1 0 1760 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_105
timestamp 1681620392
transform 1 0 1768 0 -1 570
box -8 -3 46 105
use BUFX2  BUFX2_41
timestamp 1681620392
transform 1 0 1808 0 -1 570
box -5 -3 28 105
use FILL  FILL_1283
timestamp 1681620392
transform 1 0 1832 0 -1 570
box -8 -3 16 105
use BUFX2  BUFX2_42
timestamp 1681620392
transform -1 0 1864 0 -1 570
box -5 -3 28 105
use BUFX2  BUFX2_43
timestamp 1681620392
transform 1 0 1864 0 -1 570
box -5 -3 28 105
use BUFX2  BUFX2_44
timestamp 1681620392
transform 1 0 1888 0 -1 570
box -5 -3 28 105
use OAI21X1  OAI21X1_282
timestamp 1681620392
transform 1 0 1912 0 -1 570
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_271
timestamp 1681620392
transform 1 0 1944 0 -1 570
box -8 -3 104 105
use OAI22X1  OAI22X1_106
timestamp 1681620392
transform -1 0 2080 0 -1 570
box -8 -3 46 105
use M3_M2  M3_M2_4264
timestamp 1681620392
transform 1 0 2092 0 1 475
box -3 -3 3 3
use INVX2  INVX2_328
timestamp 1681620392
transform 1 0 2080 0 -1 570
box -9 -3 26 105
use OAI22X1  OAI22X1_107
timestamp 1681620392
transform -1 0 2136 0 -1 570
box -8 -3 46 105
use M3_M2  M3_M2_4265
timestamp 1681620392
transform 1 0 2220 0 1 475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_272
timestamp 1681620392
transform 1 0 2136 0 -1 570
box -8 -3 104 105
use INVX2  INVX2_329
timestamp 1681620392
transform 1 0 2232 0 -1 570
box -9 -3 26 105
use OAI21X1  OAI21X1_283
timestamp 1681620392
transform 1 0 2248 0 -1 570
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_273
timestamp 1681620392
transform 1 0 2280 0 -1 570
box -8 -3 104 105
use NAND2X1  NAND2X1_287
timestamp 1681620392
transform 1 0 2376 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_288
timestamp 1681620392
transform 1 0 2400 0 -1 570
box -8 -3 32 105
use OAI21X1  OAI21X1_284
timestamp 1681620392
transform -1 0 2456 0 -1 570
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_274
timestamp 1681620392
transform 1 0 2456 0 -1 570
box -8 -3 104 105
use FILL  FILL_1284
timestamp 1681620392
transform 1 0 2552 0 -1 570
box -8 -3 16 105
use FILL  FILL_1285
timestamp 1681620392
transform 1 0 2560 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_275
timestamp 1681620392
transform 1 0 2568 0 -1 570
box -8 -3 104 105
use FILL  FILL_1286
timestamp 1681620392
transform 1 0 2664 0 -1 570
box -8 -3 16 105
use FILL  FILL_1287
timestamp 1681620392
transform 1 0 2672 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_44
timestamp 1681620392
transform -1 0 2720 0 -1 570
box -8 -3 46 105
use FILL  FILL_1288
timestamp 1681620392
transform 1 0 2720 0 -1 570
box -8 -3 16 105
use FILL  FILL_1289
timestamp 1681620392
transform 1 0 2728 0 -1 570
box -8 -3 16 105
use FILL  FILL_1290
timestamp 1681620392
transform 1 0 2736 0 -1 570
box -8 -3 16 105
use FILL  FILL_1291
timestamp 1681620392
transform 1 0 2744 0 -1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_285
timestamp 1681620392
transform 1 0 2752 0 -1 570
box -8 -3 34 105
use FILL  FILL_1292
timestamp 1681620392
transform 1 0 2784 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_330
timestamp 1681620392
transform 1 0 2792 0 -1 570
box -9 -3 26 105
use FILL  FILL_1293
timestamp 1681620392
transform 1 0 2808 0 -1 570
box -8 -3 16 105
use FILL  FILL_1294
timestamp 1681620392
transform 1 0 2816 0 -1 570
box -8 -3 16 105
use FILL  FILL_1295
timestamp 1681620392
transform 1 0 2824 0 -1 570
box -8 -3 16 105
use FILL  FILL_1296
timestamp 1681620392
transform 1 0 2832 0 -1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_94
timestamp 1681620392
transform -1 0 2864 0 -1 570
box -8 -3 32 105
use FILL  FILL_1297
timestamp 1681620392
transform 1 0 2864 0 -1 570
box -8 -3 16 105
use FILL  FILL_1298
timestamp 1681620392
transform 1 0 2872 0 -1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_286
timestamp 1681620392
transform 1 0 2880 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_287
timestamp 1681620392
transform -1 0 2944 0 -1 570
box -8 -3 34 105
use INVX2  INVX2_331
timestamp 1681620392
transform -1 0 2960 0 -1 570
box -9 -3 26 105
use FILL  FILL_1299
timestamp 1681620392
transform 1 0 2960 0 -1 570
box -8 -3 16 105
use FILL  FILL_1301
timestamp 1681620392
transform 1 0 2968 0 -1 570
box -8 -3 16 105
use FILL  FILL_1303
timestamp 1681620392
transform 1 0 2976 0 -1 570
box -8 -3 16 105
use FILL  FILL_1305
timestamp 1681620392
transform 1 0 2984 0 -1 570
box -8 -3 16 105
use FILL  FILL_1306
timestamp 1681620392
transform 1 0 2992 0 -1 570
box -8 -3 16 105
use FILL  FILL_1307
timestamp 1681620392
transform 1 0 3000 0 -1 570
box -8 -3 16 105
use FILL  FILL_1309
timestamp 1681620392
transform 1 0 3008 0 -1 570
box -8 -3 16 105
use Project_Top_VIA0  Project_Top_VIA0_51
timestamp 1681620392
transform 1 0 3067 0 1 470
box -10 -3 10 3
use M3_M2  M3_M2_4303
timestamp 1681620392
transform 1 0 156 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4304
timestamp 1681620392
transform 1 0 188 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4325
timestamp 1681620392
transform 1 0 124 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_4960
timestamp 1681620392
transform 1 0 132 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4961
timestamp 1681620392
transform 1 0 156 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4326
timestamp 1681620392
transform 1 0 164 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_4962
timestamp 1681620392
transform 1 0 172 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4963
timestamp 1681620392
transform 1 0 188 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4964
timestamp 1681620392
transform 1 0 196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5034
timestamp 1681620392
transform 1 0 124 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5035
timestamp 1681620392
transform 1 0 140 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5036
timestamp 1681620392
transform 1 0 156 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5037
timestamp 1681620392
transform 1 0 164 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5038
timestamp 1681620392
transform 1 0 180 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4362
timestamp 1681620392
transform 1 0 156 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4363
timestamp 1681620392
transform 1 0 196 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_5039
timestamp 1681620392
transform 1 0 212 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5040
timestamp 1681620392
transform 1 0 220 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4364
timestamp 1681620392
transform 1 0 212 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_4965
timestamp 1681620392
transform 1 0 236 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4365
timestamp 1681620392
transform 1 0 236 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_5041
timestamp 1681620392
transform 1 0 260 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4366
timestamp 1681620392
transform 1 0 260 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4281
timestamp 1681620392
transform 1 0 284 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4305
timestamp 1681620392
transform 1 0 276 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_4966
timestamp 1681620392
transform 1 0 276 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4967
timestamp 1681620392
transform 1 0 292 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4968
timestamp 1681620392
transform 1 0 300 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5042
timestamp 1681620392
transform 1 0 284 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4367
timestamp 1681620392
transform 1 0 300 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4327
timestamp 1681620392
transform 1 0 324 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4306
timestamp 1681620392
transform 1 0 340 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_4969
timestamp 1681620392
transform 1 0 340 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5043
timestamp 1681620392
transform 1 0 324 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5044
timestamp 1681620392
transform 1 0 332 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5121
timestamp 1681620392
transform 1 0 316 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_4392
timestamp 1681620392
transform 1 0 316 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_4928
timestamp 1681620392
transform 1 0 380 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4970
timestamp 1681620392
transform 1 0 380 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5045
timestamp 1681620392
transform 1 0 388 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4368
timestamp 1681620392
transform 1 0 380 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4393
timestamp 1681620392
transform 1 0 388 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_4929
timestamp 1681620392
transform 1 0 412 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5046
timestamp 1681620392
transform 1 0 404 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4369
timestamp 1681620392
transform 1 0 404 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4282
timestamp 1681620392
transform 1 0 428 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4307
timestamp 1681620392
transform 1 0 428 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_4971
timestamp 1681620392
transform 1 0 428 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4283
timestamp 1681620392
transform 1 0 460 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_5047
timestamp 1681620392
transform 1 0 452 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5048
timestamp 1681620392
transform 1 0 468 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4284
timestamp 1681620392
transform 1 0 484 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_4930
timestamp 1681620392
transform 1 0 484 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_4285
timestamp 1681620392
transform 1 0 508 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_4923
timestamp 1681620392
transform 1 0 532 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_4931
timestamp 1681620392
transform 1 0 516 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_4328
timestamp 1681620392
transform 1 0 484 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_4972
timestamp 1681620392
transform 1 0 492 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4329
timestamp 1681620392
transform 1 0 500 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_4973
timestamp 1681620392
transform 1 0 508 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4330
timestamp 1681620392
transform 1 0 516 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4286
timestamp 1681620392
transform 1 0 548 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4272
timestamp 1681620392
transform 1 0 580 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_4924
timestamp 1681620392
transform 1 0 564 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_4932
timestamp 1681620392
transform 1 0 540 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4933
timestamp 1681620392
transform 1 0 548 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4974
timestamp 1681620392
transform 1 0 524 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4394
timestamp 1681620392
transform 1 0 476 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_5049
timestamp 1681620392
transform 1 0 508 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4370
timestamp 1681620392
transform 1 0 532 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4395
timestamp 1681620392
transform 1 0 508 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4308
timestamp 1681620392
transform 1 0 556 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4287
timestamp 1681620392
transform 1 0 588 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_4925
timestamp 1681620392
transform 1 0 596 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_4934
timestamp 1681620392
transform 1 0 572 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4935
timestamp 1681620392
transform 1 0 580 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4975
timestamp 1681620392
transform 1 0 556 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4396
timestamp 1681620392
transform 1 0 540 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4331
timestamp 1681620392
transform 1 0 572 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_4936
timestamp 1681620392
transform 1 0 604 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4976
timestamp 1681620392
transform 1 0 588 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4332
timestamp 1681620392
transform 1 0 612 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_5050
timestamp 1681620392
transform 1 0 612 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4309
timestamp 1681620392
transform 1 0 628 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4273
timestamp 1681620392
transform 1 0 668 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_4937
timestamp 1681620392
transform 1 0 660 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_4274
timestamp 1681620392
transform 1 0 700 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_4926
timestamp 1681620392
transform 1 0 708 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_4938
timestamp 1681620392
transform 1 0 692 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4977
timestamp 1681620392
transform 1 0 668 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4978
timestamp 1681620392
transform 1 0 676 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4288
timestamp 1681620392
transform 1 0 716 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4275
timestamp 1681620392
transform 1 0 756 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_4939
timestamp 1681620392
transform 1 0 716 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_4310
timestamp 1681620392
transform 1 0 740 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4289
timestamp 1681620392
transform 1 0 764 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_4940
timestamp 1681620392
transform 1 0 748 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4979
timestamp 1681620392
transform 1 0 700 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4980
timestamp 1681620392
transform 1 0 724 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5051
timestamp 1681620392
transform 1 0 684 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5052
timestamp 1681620392
transform 1 0 724 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4981
timestamp 1681620392
transform 1 0 764 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4333
timestamp 1681620392
transform 1 0 780 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4290
timestamp 1681620392
transform 1 0 836 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4311
timestamp 1681620392
transform 1 0 884 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_4941
timestamp 1681620392
transform 1 0 892 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4982
timestamp 1681620392
transform 1 0 788 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4983
timestamp 1681620392
transform 1 0 828 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4984
timestamp 1681620392
transform 1 0 884 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4334
timestamp 1681620392
transform 1 0 892 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4266
timestamp 1681620392
transform 1 0 916 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_4291
timestamp 1681620392
transform 1 0 908 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_4985
timestamp 1681620392
transform 1 0 900 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5053
timestamp 1681620392
transform 1 0 748 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5054
timestamp 1681620392
transform 1 0 756 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5055
timestamp 1681620392
transform 1 0 772 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5056
timestamp 1681620392
transform 1 0 788 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5057
timestamp 1681620392
transform 1 0 804 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4371
timestamp 1681620392
transform 1 0 772 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4372
timestamp 1681620392
transform 1 0 828 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4397
timestamp 1681620392
transform 1 0 756 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4398
timestamp 1681620392
transform 1 0 788 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4399
timestamp 1681620392
transform 1 0 844 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4267
timestamp 1681620392
transform 1 0 1028 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_4312
timestamp 1681620392
transform 1 0 1028 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4276
timestamp 1681620392
transform 1 0 1068 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_4942
timestamp 1681620392
transform 1 0 1068 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4986
timestamp 1681620392
transform 1 0 924 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4987
timestamp 1681620392
transform 1 0 964 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4988
timestamp 1681620392
transform 1 0 1020 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4989
timestamp 1681620392
transform 1 0 1036 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4990
timestamp 1681620392
transform 1 0 1052 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5058
timestamp 1681620392
transform 1 0 908 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5059
timestamp 1681620392
transform 1 0 916 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4313
timestamp 1681620392
transform 1 0 1092 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4314
timestamp 1681620392
transform 1 0 1132 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_4991
timestamp 1681620392
transform 1 0 1084 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5060
timestamp 1681620392
transform 1 0 940 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5061
timestamp 1681620392
transform 1 0 1028 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5062
timestamp 1681620392
transform 1 0 1044 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5063
timestamp 1681620392
transform 1 0 1060 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5064
timestamp 1681620392
transform 1 0 1068 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4400
timestamp 1681620392
transform 1 0 940 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4401
timestamp 1681620392
transform 1 0 980 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4353
timestamp 1681620392
transform 1 0 1084 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_4992
timestamp 1681620392
transform 1 0 1132 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4993
timestamp 1681620392
transform 1 0 1188 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5065
timestamp 1681620392
transform 1 0 1092 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5066
timestamp 1681620392
transform 1 0 1108 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4373
timestamp 1681620392
transform 1 0 1068 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4354
timestamp 1681620392
transform 1 0 1180 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_5067
timestamp 1681620392
transform 1 0 1196 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4374
timestamp 1681620392
transform 1 0 1132 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_4994
timestamp 1681620392
transform 1 0 1220 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4995
timestamp 1681620392
transform 1 0 1244 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4335
timestamp 1681620392
transform 1 0 1252 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4336
timestamp 1681620392
transform 1 0 1268 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_4996
timestamp 1681620392
transform 1 0 1284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4997
timestamp 1681620392
transform 1 0 1332 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4998
timestamp 1681620392
transform 1 0 1380 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5068
timestamp 1681620392
transform 1 0 1236 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5069
timestamp 1681620392
transform 1 0 1260 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5070
timestamp 1681620392
transform 1 0 1268 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4375
timestamp 1681620392
transform 1 0 1260 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_5071
timestamp 1681620392
transform 1 0 1300 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5072
timestamp 1681620392
transform 1 0 1388 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5073
timestamp 1681620392
transform 1 0 1396 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4376
timestamp 1681620392
transform 1 0 1300 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_4927
timestamp 1681620392
transform 1 0 1444 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_4943
timestamp 1681620392
transform 1 0 1428 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_4337
timestamp 1681620392
transform 1 0 1428 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_4944
timestamp 1681620392
transform 1 0 1460 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5074
timestamp 1681620392
transform 1 0 1420 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5075
timestamp 1681620392
transform 1 0 1436 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5076
timestamp 1681620392
transform 1 0 1460 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4292
timestamp 1681620392
transform 1 0 1476 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_4945
timestamp 1681620392
transform 1 0 1476 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4946
timestamp 1681620392
transform 1 0 1484 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4999
timestamp 1681620392
transform 1 0 1476 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4338
timestamp 1681620392
transform 1 0 1484 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4277
timestamp 1681620392
transform 1 0 1532 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_4293
timestamp 1681620392
transform 1 0 1524 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_4947
timestamp 1681620392
transform 1 0 1508 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5000
timestamp 1681620392
transform 1 0 1500 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4402
timestamp 1681620392
transform 1 0 1476 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4339
timestamp 1681620392
transform 1 0 1508 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_5077
timestamp 1681620392
transform 1 0 1516 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4948
timestamp 1681620392
transform 1 0 1532 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_4315
timestamp 1681620392
transform 1 0 1540 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4340
timestamp 1681620392
transform 1 0 1532 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4294
timestamp 1681620392
transform 1 0 1572 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_5001
timestamp 1681620392
transform 1 0 1540 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5002
timestamp 1681620392
transform 1 0 1548 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5078
timestamp 1681620392
transform 1 0 1540 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5079
timestamp 1681620392
transform 1 0 1564 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4949
timestamp 1681620392
transform 1 0 1572 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_4316
timestamp 1681620392
transform 1 0 1588 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_5003
timestamp 1681620392
transform 1 0 1588 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4341
timestamp 1681620392
transform 1 0 1596 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4278
timestamp 1681620392
transform 1 0 1628 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_4295
timestamp 1681620392
transform 1 0 1636 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_4950
timestamp 1681620392
transform 1 0 1628 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4951
timestamp 1681620392
transform 1 0 1636 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_4342
timestamp 1681620392
transform 1 0 1628 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_5004
timestamp 1681620392
transform 1 0 1636 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5080
timestamp 1681620392
transform 1 0 1596 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5081
timestamp 1681620392
transform 1 0 1604 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5082
timestamp 1681620392
transform 1 0 1612 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4355
timestamp 1681620392
transform 1 0 1620 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_5083
timestamp 1681620392
transform 1 0 1628 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5005
timestamp 1681620392
transform 1 0 1676 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5084
timestamp 1681620392
transform 1 0 1660 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4356
timestamp 1681620392
transform 1 0 1668 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_4317
timestamp 1681620392
transform 1 0 1748 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_5006
timestamp 1681620392
transform 1 0 1692 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5007
timestamp 1681620392
transform 1 0 1748 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4343
timestamp 1681620392
transform 1 0 1772 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_5085
timestamp 1681620392
transform 1 0 1772 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4377
timestamp 1681620392
transform 1 0 1740 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4403
timestamp 1681620392
transform 1 0 1772 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4318
timestamp 1681620392
transform 1 0 1788 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_5086
timestamp 1681620392
transform 1 0 1788 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4378
timestamp 1681620392
transform 1 0 1788 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4296
timestamp 1681620392
transform 1 0 1796 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4344
timestamp 1681620392
transform 1 0 1820 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_5087
timestamp 1681620392
transform 1 0 1820 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4268
timestamp 1681620392
transform 1 0 1868 0 1 455
box -3 -3 3 3
use M2_M1  M2_M1_5008
timestamp 1681620392
transform 1 0 1852 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5009
timestamp 1681620392
transform 1 0 1868 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5088
timestamp 1681620392
transform 1 0 1844 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4357
timestamp 1681620392
transform 1 0 1852 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_5089
timestamp 1681620392
transform 1 0 1860 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5090
timestamp 1681620392
transform 1 0 1876 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4379
timestamp 1681620392
transform 1 0 1844 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4380
timestamp 1681620392
transform 1 0 1884 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4279
timestamp 1681620392
transform 1 0 1972 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_4297
timestamp 1681620392
transform 1 0 1996 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4319
timestamp 1681620392
transform 1 0 2036 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_5010
timestamp 1681620392
transform 1 0 1996 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4345
timestamp 1681620392
transform 1 0 2028 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_5011
timestamp 1681620392
transform 1 0 2036 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5091
timestamp 1681620392
transform 1 0 1948 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4404
timestamp 1681620392
transform 1 0 1988 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4269
timestamp 1681620392
transform 1 0 2052 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_4298
timestamp 1681620392
transform 1 0 2060 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4320
timestamp 1681620392
transform 1 0 2084 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_5012
timestamp 1681620392
transform 1 0 2052 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4346
timestamp 1681620392
transform 1 0 2060 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_5013
timestamp 1681620392
transform 1 0 2068 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4280
timestamp 1681620392
transform 1 0 2108 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_4299
timestamp 1681620392
transform 1 0 2108 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_4952
timestamp 1681620392
transform 1 0 2108 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5014
timestamp 1681620392
transform 1 0 2092 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5092
timestamp 1681620392
transform 1 0 2036 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5093
timestamp 1681620392
transform 1 0 2044 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5094
timestamp 1681620392
transform 1 0 2060 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5095
timestamp 1681620392
transform 1 0 2076 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5096
timestamp 1681620392
transform 1 0 2084 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4358
timestamp 1681620392
transform 1 0 2092 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_5015
timestamp 1681620392
transform 1 0 2148 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5097
timestamp 1681620392
transform 1 0 2108 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5098
timestamp 1681620392
transform 1 0 2124 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4381
timestamp 1681620392
transform 1 0 2108 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4382
timestamp 1681620392
transform 1 0 2148 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_5016
timestamp 1681620392
transform 1 0 2212 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5017
timestamp 1681620392
transform 1 0 2220 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5099
timestamp 1681620392
transform 1 0 2220 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4383
timestamp 1681620392
transform 1 0 2212 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4300
timestamp 1681620392
transform 1 0 2284 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_4953
timestamp 1681620392
transform 1 0 2268 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_4321
timestamp 1681620392
transform 1 0 2276 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4347
timestamp 1681620392
transform 1 0 2268 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_4954
timestamp 1681620392
transform 1 0 2292 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_4322
timestamp 1681620392
transform 1 0 2308 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_5018
timestamp 1681620392
transform 1 0 2284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5100
timestamp 1681620392
transform 1 0 2244 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5101
timestamp 1681620392
transform 1 0 2252 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5102
timestamp 1681620392
transform 1 0 2268 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4384
timestamp 1681620392
transform 1 0 2268 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4348
timestamp 1681620392
transform 1 0 2292 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_5019
timestamp 1681620392
transform 1 0 2308 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4270
timestamp 1681620392
transform 1 0 2388 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_4271
timestamp 1681620392
transform 1 0 2412 0 1 455
box -3 -3 3 3
use M2_M1  M2_M1_5020
timestamp 1681620392
transform 1 0 2356 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5021
timestamp 1681620392
transform 1 0 2412 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5103
timestamp 1681620392
transform 1 0 2316 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5104
timestamp 1681620392
transform 1 0 2332 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4385
timestamp 1681620392
transform 1 0 2316 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_5105
timestamp 1681620392
transform 1 0 2420 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4386
timestamp 1681620392
transform 1 0 2412 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4405
timestamp 1681620392
transform 1 0 2420 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_4955
timestamp 1681620392
transform 1 0 2444 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_4301
timestamp 1681620392
transform 1 0 2460 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_5022
timestamp 1681620392
transform 1 0 2460 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4302
timestamp 1681620392
transform 1 0 2564 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_4956
timestamp 1681620392
transform 1 0 2564 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5023
timestamp 1681620392
transform 1 0 2500 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5024
timestamp 1681620392
transform 1 0 2556 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5106
timestamp 1681620392
transform 1 0 2476 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5025
timestamp 1681620392
transform 1 0 2596 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5107
timestamp 1681620392
transform 1 0 2580 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5108
timestamp 1681620392
transform 1 0 2628 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4387
timestamp 1681620392
transform 1 0 2644 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_5026
timestamp 1681620392
transform 1 0 2692 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5109
timestamp 1681620392
transform 1 0 2668 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5110
timestamp 1681620392
transform 1 0 2684 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4406
timestamp 1681620392
transform 1 0 2676 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4349
timestamp 1681620392
transform 1 0 2716 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_5027
timestamp 1681620392
transform 1 0 2724 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5028
timestamp 1681620392
transform 1 0 2740 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5111
timestamp 1681620392
transform 1 0 2708 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4350
timestamp 1681620392
transform 1 0 2748 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_5029
timestamp 1681620392
transform 1 0 2756 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5112
timestamp 1681620392
transform 1 0 2732 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5113
timestamp 1681620392
transform 1 0 2748 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5114
timestamp 1681620392
transform 1 0 2756 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4388
timestamp 1681620392
transform 1 0 2732 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4407
timestamp 1681620392
transform 1 0 2740 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4359
timestamp 1681620392
transform 1 0 2764 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_4323
timestamp 1681620392
transform 1 0 2788 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4324
timestamp 1681620392
transform 1 0 2820 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4351
timestamp 1681620392
transform 1 0 2820 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_5115
timestamp 1681620392
transform 1 0 2820 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4957
timestamp 1681620392
transform 1 0 2860 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5030
timestamp 1681620392
transform 1 0 2836 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5031
timestamp 1681620392
transform 1 0 2844 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_4360
timestamp 1681620392
transform 1 0 2844 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_4352
timestamp 1681620392
transform 1 0 2868 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_5032
timestamp 1681620392
transform 1 0 2884 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5116
timestamp 1681620392
transform 1 0 2884 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4408
timestamp 1681620392
transform 1 0 2884 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_5117
timestamp 1681620392
transform 1 0 2900 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5118
timestamp 1681620392
transform 1 0 2908 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4958
timestamp 1681620392
transform 1 0 2924 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5033
timestamp 1681620392
transform 1 0 2932 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5119
timestamp 1681620392
transform 1 0 2924 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_4361
timestamp 1681620392
transform 1 0 2932 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_4389
timestamp 1681620392
transform 1 0 2916 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4390
timestamp 1681620392
transform 1 0 2932 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_5120
timestamp 1681620392
transform 1 0 2956 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4959
timestamp 1681620392
transform 1 0 2964 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_4391
timestamp 1681620392
transform 1 0 2964 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4409
timestamp 1681620392
transform 1 0 2956 0 1 385
box -3 -3 3 3
use Project_Top_VIA0  Project_Top_VIA0_52
timestamp 1681620392
transform 1 0 48 0 1 370
box -10 -3 10 3
use FILL  FILL_1310
timestamp 1681620392
transform 1 0 72 0 1 370
box -8 -3 16 105
use FILL  FILL_1311
timestamp 1681620392
transform 1 0 80 0 1 370
box -8 -3 16 105
use FILL  FILL_1312
timestamp 1681620392
transform 1 0 88 0 1 370
box -8 -3 16 105
use FILL  FILL_1313
timestamp 1681620392
transform 1 0 96 0 1 370
box -8 -3 16 105
use FILL  FILL_1314
timestamp 1681620392
transform 1 0 104 0 1 370
box -8 -3 16 105
use FILL  FILL_1315
timestamp 1681620392
transform 1 0 112 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_4410
timestamp 1681620392
transform 1 0 132 0 1 375
box -3 -3 3 3
use OAI22X1  OAI22X1_108
timestamp 1681620392
transform -1 0 160 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_109
timestamp 1681620392
transform -1 0 200 0 1 370
box -8 -3 46 105
use M3_M2  M3_M2_4411
timestamp 1681620392
transform 1 0 212 0 1 375
box -3 -3 3 3
use FILL  FILL_1316
timestamp 1681620392
transform 1 0 200 0 1 370
box -8 -3 16 105
use FILL  FILL_1317
timestamp 1681620392
transform 1 0 208 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_4412
timestamp 1681620392
transform 1 0 244 0 1 375
box -3 -3 3 3
use INVX2  INVX2_333
timestamp 1681620392
transform 1 0 216 0 1 370
box -9 -3 26 105
use INVX2  INVX2_334
timestamp 1681620392
transform -1 0 248 0 1 370
box -9 -3 26 105
use FILL  FILL_1318
timestamp 1681620392
transform 1 0 248 0 1 370
box -8 -3 16 105
use FILL  FILL_1319
timestamp 1681620392
transform 1 0 256 0 1 370
box -8 -3 16 105
use FILL  FILL_1320
timestamp 1681620392
transform 1 0 264 0 1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_95
timestamp 1681620392
transform 1 0 272 0 1 370
box -8 -3 32 105
use M3_M2  M3_M2_4413
timestamp 1681620392
transform 1 0 324 0 1 375
box -3 -3 3 3
use NOR2X1  NOR2X1_96
timestamp 1681620392
transform -1 0 320 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_97
timestamp 1681620392
transform 1 0 320 0 1 370
box -8 -3 32 105
use FILL  FILL_1321
timestamp 1681620392
transform 1 0 344 0 1 370
box -8 -3 16 105
use FILL  FILL_1322
timestamp 1681620392
transform 1 0 352 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_289
timestamp 1681620392
transform 1 0 360 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_290
timestamp 1681620392
transform 1 0 384 0 1 370
box -8 -3 32 105
use FILL  FILL_1323
timestamp 1681620392
transform 1 0 408 0 1 370
box -8 -3 16 105
use FILL  FILL_1324
timestamp 1681620392
transform 1 0 416 0 1 370
box -8 -3 16 105
use INVX2  INVX2_335
timestamp 1681620392
transform 1 0 424 0 1 370
box -9 -3 26 105
use FILL  FILL_1325
timestamp 1681620392
transform 1 0 440 0 1 370
box -8 -3 16 105
use FILL  FILL_1326
timestamp 1681620392
transform 1 0 448 0 1 370
box -8 -3 16 105
use FILL  FILL_1327
timestamp 1681620392
transform 1 0 456 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_291
timestamp 1681620392
transform 1 0 464 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_292
timestamp 1681620392
transform -1 0 512 0 1 370
box -8 -3 32 105
use NAND3X1  NAND3X1_101
timestamp 1681620392
transform 1 0 512 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_102
timestamp 1681620392
transform 1 0 544 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_103
timestamp 1681620392
transform 1 0 576 0 1 370
box -8 -3 40 105
use FILL  FILL_1328
timestamp 1681620392
transform 1 0 608 0 1 370
box -8 -3 16 105
use FILL  FILL_1329
timestamp 1681620392
transform 1 0 616 0 1 370
box -8 -3 16 105
use FILL  FILL_1330
timestamp 1681620392
transform 1 0 624 0 1 370
box -8 -3 16 105
use FILL  FILL_1331
timestamp 1681620392
transform 1 0 632 0 1 370
box -8 -3 16 105
use INVX2  INVX2_336
timestamp 1681620392
transform 1 0 640 0 1 370
box -9 -3 26 105
use FILL  FILL_1332
timestamp 1681620392
transform 1 0 656 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_293
timestamp 1681620392
transform -1 0 688 0 1 370
box -8 -3 32 105
use NAND3X1  NAND3X1_104
timestamp 1681620392
transform 1 0 688 0 1 370
box -8 -3 40 105
use M3_M2  M3_M2_4414
timestamp 1681620392
transform 1 0 740 0 1 375
box -3 -3 3 3
use OAI21X1  OAI21X1_288
timestamp 1681620392
transform 1 0 720 0 1 370
box -8 -3 34 105
use M3_M2  M3_M2_4415
timestamp 1681620392
transform 1 0 796 0 1 375
box -3 -3 3 3
use OAI22X1  OAI22X1_110
timestamp 1681620392
transform -1 0 792 0 1 370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_276
timestamp 1681620392
transform 1 0 792 0 1 370
box -8 -3 104 105
use NAND2X1  NAND2X1_294
timestamp 1681620392
transform -1 0 912 0 1 370
box -8 -3 32 105
use INVX2  INVX2_337
timestamp 1681620392
transform 1 0 912 0 1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_277
timestamp 1681620392
transform 1 0 928 0 1 370
box -8 -3 104 105
use OAI22X1  OAI22X1_111
timestamp 1681620392
transform 1 0 1024 0 1 370
box -8 -3 46 105
use M3_M2  M3_M2_4416
timestamp 1681620392
transform 1 0 1108 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4417
timestamp 1681620392
transform 1 0 1164 0 1 375
box -3 -3 3 3
use OAI21X1  OAI21X1_289
timestamp 1681620392
transform -1 0 1096 0 1 370
box -8 -3 34 105
use M3_M2  M3_M2_4418
timestamp 1681620392
transform 1 0 1196 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_278
timestamp 1681620392
transform 1 0 1096 0 1 370
box -8 -3 104 105
use BUFX2  BUFX2_45
timestamp 1681620392
transform -1 0 1216 0 1 370
box -5 -3 28 105
use BUFX2  BUFX2_46
timestamp 1681620392
transform 1 0 1216 0 1 370
box -5 -3 28 105
use BUFX2  BUFX2_47
timestamp 1681620392
transform 1 0 1240 0 1 370
box -5 -3 28 105
use M3_M2  M3_M2_4419
timestamp 1681620392
transform 1 0 1284 0 1 375
box -3 -3 3 3
use BUFX2  BUFX2_48
timestamp 1681620392
transform -1 0 1288 0 1 370
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_279
timestamp 1681620392
transform 1 0 1288 0 1 370
box -8 -3 104 105
use NOR2X1  NOR2X1_98
timestamp 1681620392
transform -1 0 1408 0 1 370
box -8 -3 32 105
use INVX2  INVX2_338
timestamp 1681620392
transform -1 0 1424 0 1 370
box -9 -3 26 105
use NAND3X1  NAND3X1_105
timestamp 1681620392
transform 1 0 1424 0 1 370
box -8 -3 40 105
use NAND2X1  NAND2X1_296
timestamp 1681620392
transform 1 0 1456 0 1 370
box -8 -3 32 105
use NAND3X1  NAND3X1_114
timestamp 1681620392
transform -1 0 1512 0 1 370
box -8 -3 40 105
use NAND2X1  NAND2X1_297
timestamp 1681620392
transform 1 0 1512 0 1 370
box -8 -3 32 105
use OAI21X1  OAI21X1_292
timestamp 1681620392
transform 1 0 1536 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_293
timestamp 1681620392
transform -1 0 1600 0 1 370
box -8 -3 34 105
use FILL  FILL_1345
timestamp 1681620392
transform 1 0 1600 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_299
timestamp 1681620392
transform 1 0 1608 0 1 370
box -8 -3 32 105
use OAI21X1  OAI21X1_294
timestamp 1681620392
transform -1 0 1664 0 1 370
box -8 -3 34 105
use FILL  FILL_1346
timestamp 1681620392
transform 1 0 1664 0 1 370
box -8 -3 16 105
use FILL  FILL_1347
timestamp 1681620392
transform 1 0 1672 0 1 370
box -8 -3 16 105
use FILL  FILL_1350
timestamp 1681620392
transform 1 0 1680 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_4420
timestamp 1681620392
transform 1 0 1716 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_285
timestamp 1681620392
transform -1 0 1784 0 1 370
box -8 -3 104 105
use FILL  FILL_1351
timestamp 1681620392
transform 1 0 1784 0 1 370
box -8 -3 16 105
use FILL  FILL_1352
timestamp 1681620392
transform 1 0 1792 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_4421
timestamp 1681620392
transform 1 0 1812 0 1 375
box -3 -3 3 3
use INVX2  INVX2_350
timestamp 1681620392
transform 1 0 1800 0 1 370
box -9 -3 26 105
use FILL  FILL_1353
timestamp 1681620392
transform 1 0 1816 0 1 370
box -8 -3 16 105
use FILL  FILL_1354
timestamp 1681620392
transform 1 0 1824 0 1 370
box -8 -3 16 105
use FILL  FILL_1355
timestamp 1681620392
transform 1 0 1832 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_116
timestamp 1681620392
transform 1 0 1840 0 1 370
box -8 -3 46 105
use FILL  FILL_1361
timestamp 1681620392
transform 1 0 1880 0 1 370
box -8 -3 16 105
use FILL  FILL_1362
timestamp 1681620392
transform 1 0 1888 0 1 370
box -8 -3 16 105
use FILL  FILL_1365
timestamp 1681620392
transform 1 0 1896 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_4422
timestamp 1681620392
transform 1 0 1916 0 1 375
box -3 -3 3 3
use FILL  FILL_1366
timestamp 1681620392
transform 1 0 1904 0 1 370
box -8 -3 16 105
use FILL  FILL_1367
timestamp 1681620392
transform 1 0 1912 0 1 370
box -8 -3 16 105
use FILL  FILL_1368
timestamp 1681620392
transform 1 0 1920 0 1 370
box -8 -3 16 105
use FILL  FILL_1369
timestamp 1681620392
transform 1 0 1928 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_287
timestamp 1681620392
transform 1 0 1936 0 1 370
box -8 -3 104 105
use FILL  FILL_1370
timestamp 1681620392
transform 1 0 2032 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_4423
timestamp 1681620392
transform 1 0 2084 0 1 375
box -3 -3 3 3
use OAI22X1  OAI22X1_118
timestamp 1681620392
transform -1 0 2080 0 1 370
box -8 -3 46 105
use M3_M2  M3_M2_4424
timestamp 1681620392
transform 1 0 2180 0 1 375
box -3 -3 3 3
use OAI21X1  OAI21X1_295
timestamp 1681620392
transform 1 0 2080 0 1 370
box -8 -3 34 105
use M3_M2  M3_M2_4425
timestamp 1681620392
transform 1 0 2204 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_288
timestamp 1681620392
transform 1 0 2112 0 1 370
box -8 -3 104 105
use FILL  FILL_1371
timestamp 1681620392
transform 1 0 2208 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_296
timestamp 1681620392
transform 1 0 2216 0 1 370
box -8 -3 34 105
use NAND2X1  NAND2X1_302
timestamp 1681620392
transform 1 0 2248 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_303
timestamp 1681620392
transform 1 0 2272 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_304
timestamp 1681620392
transform -1 0 2320 0 1 370
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_291
timestamp 1681620392
transform 1 0 2320 0 1 370
box -8 -3 104 105
use FILL  FILL_1387
timestamp 1681620392
transform 1 0 2416 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_306
timestamp 1681620392
transform 1 0 2424 0 1 370
box -8 -3 32 105
use FILL  FILL_1388
timestamp 1681620392
transform 1 0 2448 0 1 370
box -8 -3 16 105
use FILL  FILL_1389
timestamp 1681620392
transform 1 0 2456 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_4426
timestamp 1681620392
transform 1 0 2532 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4427
timestamp 1681620392
transform 1 0 2556 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_293
timestamp 1681620392
transform 1 0 2464 0 1 370
box -8 -3 104 105
use FILL  FILL_1390
timestamp 1681620392
transform 1 0 2560 0 1 370
box -8 -3 16 105
use FILL  FILL_1391
timestamp 1681620392
transform 1 0 2568 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_298
timestamp 1681620392
transform -1 0 2608 0 1 370
box -8 -3 34 105
use FILL  FILL_1392
timestamp 1681620392
transform 1 0 2608 0 1 370
box -8 -3 16 105
use INVX2  INVX2_352
timestamp 1681620392
transform -1 0 2632 0 1 370
box -9 -3 26 105
use FILL  FILL_1393
timestamp 1681620392
transform 1 0 2632 0 1 370
box -8 -3 16 105
use FILL  FILL_1394
timestamp 1681620392
transform 1 0 2640 0 1 370
box -8 -3 16 105
use FILL  FILL_1395
timestamp 1681620392
transform 1 0 2648 0 1 370
box -8 -3 16 105
use FILL  FILL_1400
timestamp 1681620392
transform 1 0 2656 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_120
timestamp 1681620392
transform 1 0 2664 0 1 370
box -8 -3 46 105
use FILL  FILL_1401
timestamp 1681620392
transform 1 0 2704 0 1 370
box -8 -3 16 105
use FILL  FILL_1402
timestamp 1681620392
transform 1 0 2712 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_45
timestamp 1681620392
transform -1 0 2760 0 1 370
box -8 -3 46 105
use FILL  FILL_1403
timestamp 1681620392
transform 1 0 2760 0 1 370
box -8 -3 16 105
use FILL  FILL_1407
timestamp 1681620392
transform 1 0 2768 0 1 370
box -8 -3 16 105
use FILL  FILL_1409
timestamp 1681620392
transform 1 0 2776 0 1 370
box -8 -3 16 105
use FILL  FILL_1410
timestamp 1681620392
transform 1 0 2784 0 1 370
box -8 -3 16 105
use FILL  FILL_1411
timestamp 1681620392
transform 1 0 2792 0 1 370
box -8 -3 16 105
use INVX2  INVX2_356
timestamp 1681620392
transform 1 0 2800 0 1 370
box -9 -3 26 105
use FILL  FILL_1412
timestamp 1681620392
transform 1 0 2816 0 1 370
box -8 -3 16 105
use FILL  FILL_1413
timestamp 1681620392
transform 1 0 2824 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_301
timestamp 1681620392
transform 1 0 2832 0 1 370
box -8 -3 34 105
use FILL  FILL_1414
timestamp 1681620392
transform 1 0 2864 0 1 370
box -8 -3 16 105
use FILL  FILL_1415
timestamp 1681620392
transform 1 0 2872 0 1 370
box -8 -3 16 105
use FILL  FILL_1416
timestamp 1681620392
transform 1 0 2880 0 1 370
box -8 -3 16 105
use INVX2  INVX2_357
timestamp 1681620392
transform -1 0 2904 0 1 370
box -9 -3 26 105
use M3_M2  M3_M2_4428
timestamp 1681620392
transform 1 0 2924 0 1 375
box -3 -3 3 3
use NAND2X1  NAND2X1_309
timestamp 1681620392
transform 1 0 2904 0 1 370
box -8 -3 32 105
use OAI21X1  OAI21X1_302
timestamp 1681620392
transform 1 0 2928 0 1 370
box -8 -3 34 105
use FILL  FILL_1417
timestamp 1681620392
transform 1 0 2960 0 1 370
box -8 -3 16 105
use FILL  FILL_1418
timestamp 1681620392
transform 1 0 2968 0 1 370
box -8 -3 16 105
use FILL  FILL_1421
timestamp 1681620392
transform 1 0 2976 0 1 370
box -8 -3 16 105
use FILL  FILL_1423
timestamp 1681620392
transform 1 0 2984 0 1 370
box -8 -3 16 105
use FILL  FILL_1425
timestamp 1681620392
transform 1 0 2992 0 1 370
box -8 -3 16 105
use FILL  FILL_1427
timestamp 1681620392
transform 1 0 3000 0 1 370
box -8 -3 16 105
use FILL  FILL_1429
timestamp 1681620392
transform 1 0 3008 0 1 370
box -8 -3 16 105
use Project_Top_VIA0  Project_Top_VIA0_53
timestamp 1681620392
transform 1 0 3043 0 1 370
box -10 -3 10 3
use M3_M2  M3_M2_4457
timestamp 1681620392
transform 1 0 180 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4458
timestamp 1681620392
transform 1 0 204 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_5128
timestamp 1681620392
transform 1 0 84 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4484
timestamp 1681620392
transform 1 0 164 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_5129
timestamp 1681620392
transform 1 0 180 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4485
timestamp 1681620392
transform 1 0 220 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_5198
timestamp 1681620392
transform 1 0 132 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4504
timestamp 1681620392
transform 1 0 148 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_5199
timestamp 1681620392
transform 1 0 164 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5200
timestamp 1681620392
transform 1 0 204 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5201
timestamp 1681620392
transform 1 0 260 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4527
timestamp 1681620392
transform 1 0 84 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4528
timestamp 1681620392
transform 1 0 180 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4584
timestamp 1681620392
transform 1 0 220 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_4444
timestamp 1681620392
transform 1 0 284 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_5122
timestamp 1681620392
transform 1 0 292 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_5130
timestamp 1681620392
transform 1 0 284 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4486
timestamp 1681620392
transform 1 0 292 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_5131
timestamp 1681620392
transform 1 0 300 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4459
timestamp 1681620392
transform 1 0 332 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_5132
timestamp 1681620392
transform 1 0 316 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4487
timestamp 1681620392
transform 1 0 324 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_4445
timestamp 1681620392
transform 1 0 412 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_4460
timestamp 1681620392
transform 1 0 388 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_5123
timestamp 1681620392
transform 1 0 452 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_5133
timestamp 1681620392
transform 1 0 332 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5134
timestamp 1681620392
transform 1 0 348 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5135
timestamp 1681620392
transform 1 0 364 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5202
timestamp 1681620392
transform 1 0 308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5203
timestamp 1681620392
transform 1 0 324 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4505
timestamp 1681620392
transform 1 0 332 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_5204
timestamp 1681620392
transform 1 0 340 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4506
timestamp 1681620392
transform 1 0 348 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_5205
timestamp 1681620392
transform 1 0 388 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4507
timestamp 1681620392
transform 1 0 436 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_5206
timestamp 1681620392
transform 1 0 444 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5207
timestamp 1681620392
transform 1 0 452 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4529
timestamp 1681620392
transform 1 0 452 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_5136
timestamp 1681620392
transform 1 0 484 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5208
timestamp 1681620392
transform 1 0 476 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5276
timestamp 1681620392
transform 1 0 484 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5137
timestamp 1681620392
transform 1 0 500 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5138
timestamp 1681620392
transform 1 0 540 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5209
timestamp 1681620392
transform 1 0 516 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4530
timestamp 1681620392
transform 1 0 500 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4508
timestamp 1681620392
transform 1 0 540 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_5139
timestamp 1681620392
transform 1 0 572 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5210
timestamp 1681620392
transform 1 0 548 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5211
timestamp 1681620392
transform 1 0 564 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5277
timestamp 1681620392
transform 1 0 516 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5278
timestamp 1681620392
transform 1 0 540 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5307
timestamp 1681620392
transform 1 0 500 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_4553
timestamp 1681620392
transform 1 0 516 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_4509
timestamp 1681620392
transform 1 0 572 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_4554
timestamp 1681620392
transform 1 0 548 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_4461
timestamp 1681620392
transform 1 0 604 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_5212
timestamp 1681620392
transform 1 0 604 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5279
timestamp 1681620392
transform 1 0 596 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5308
timestamp 1681620392
transform 1 0 588 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_4555
timestamp 1681620392
transform 1 0 596 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_4462
timestamp 1681620392
transform 1 0 644 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_5140
timestamp 1681620392
transform 1 0 644 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5213
timestamp 1681620392
transform 1 0 620 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4510
timestamp 1681620392
transform 1 0 636 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_5124
timestamp 1681620392
transform 1 0 676 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_5141
timestamp 1681620392
transform 1 0 668 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5142
timestamp 1681620392
transform 1 0 676 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4511
timestamp 1681620392
transform 1 0 676 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_5214
timestamp 1681620392
transform 1 0 692 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4512
timestamp 1681620392
transform 1 0 700 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_5215
timestamp 1681620392
transform 1 0 708 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5280
timestamp 1681620392
transform 1 0 636 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_4531
timestamp 1681620392
transform 1 0 668 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_5281
timestamp 1681620392
transform 1 0 700 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5216
timestamp 1681620392
transform 1 0 748 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5282
timestamp 1681620392
transform 1 0 724 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5283
timestamp 1681620392
transform 1 0 732 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_4556
timestamp 1681620392
transform 1 0 708 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_5309
timestamp 1681620392
transform 1 0 716 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_4573
timestamp 1681620392
transform 1 0 700 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4585
timestamp 1681620392
transform 1 0 716 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_4532
timestamp 1681620392
transform 1 0 740 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_5217
timestamp 1681620392
transform 1 0 772 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4513
timestamp 1681620392
transform 1 0 780 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_5284
timestamp 1681620392
transform 1 0 756 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5285
timestamp 1681620392
transform 1 0 764 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5310
timestamp 1681620392
transform 1 0 740 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_4557
timestamp 1681620392
transform 1 0 748 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_5311
timestamp 1681620392
transform 1 0 780 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_4574
timestamp 1681620392
transform 1 0 772 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4463
timestamp 1681620392
transform 1 0 804 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_5143
timestamp 1681620392
transform 1 0 796 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4586
timestamp 1681620392
transform 1 0 788 0 1 285
box -3 -3 3 3
use M2_M1  M2_M1_5144
timestamp 1681620392
transform 1 0 812 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5145
timestamp 1681620392
transform 1 0 876 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5218
timestamp 1681620392
transform 1 0 820 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5219
timestamp 1681620392
transform 1 0 836 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5220
timestamp 1681620392
transform 1 0 852 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5286
timestamp 1681620392
transform 1 0 804 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_4533
timestamp 1681620392
transform 1 0 812 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4514
timestamp 1681620392
transform 1 0 868 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_4429
timestamp 1681620392
transform 1 0 924 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_4430
timestamp 1681620392
transform 1 0 972 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_4446
timestamp 1681620392
transform 1 0 940 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_4464
timestamp 1681620392
transform 1 0 948 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4447
timestamp 1681620392
transform 1 0 980 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_5146
timestamp 1681620392
transform 1 0 900 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5147
timestamp 1681620392
transform 1 0 908 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5148
timestamp 1681620392
transform 1 0 924 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5149
timestamp 1681620392
transform 1 0 940 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5150
timestamp 1681620392
transform 1 0 948 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5151
timestamp 1681620392
transform 1 0 964 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5152
timestamp 1681620392
transform 1 0 980 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5221
timestamp 1681620392
transform 1 0 884 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5287
timestamp 1681620392
transform 1 0 844 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_4558
timestamp 1681620392
transform 1 0 820 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_4534
timestamp 1681620392
transform 1 0 860 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_5288
timestamp 1681620392
transform 1 0 868 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_4559
timestamp 1681620392
transform 1 0 852 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_5312
timestamp 1681620392
transform 1 0 860 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_4575
timestamp 1681620392
transform 1 0 836 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4587
timestamp 1681620392
transform 1 0 828 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_4588
timestamp 1681620392
transform 1 0 860 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_4515
timestamp 1681620392
transform 1 0 908 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_5222
timestamp 1681620392
transform 1 0 916 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5223
timestamp 1681620392
transform 1 0 932 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5289
timestamp 1681620392
transform 1 0 900 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_4560
timestamp 1681620392
transform 1 0 892 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_4576
timestamp 1681620392
transform 1 0 900 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_5224
timestamp 1681620392
transform 1 0 956 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4448
timestamp 1681620392
transform 1 0 1028 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_4465
timestamp 1681620392
transform 1 0 1036 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_5153
timestamp 1681620392
transform 1 0 1012 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5154
timestamp 1681620392
transform 1 0 1028 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5155
timestamp 1681620392
transform 1 0 1036 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5225
timestamp 1681620392
transform 1 0 1012 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5290
timestamp 1681620392
transform 1 0 1036 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_4561
timestamp 1681620392
transform 1 0 1036 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_4431
timestamp 1681620392
transform 1 0 1068 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_4449
timestamp 1681620392
transform 1 0 1060 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_4432
timestamp 1681620392
transform 1 0 1092 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_4450
timestamp 1681620392
transform 1 0 1092 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_4466
timestamp 1681620392
transform 1 0 1116 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_5156
timestamp 1681620392
transform 1 0 1060 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5157
timestamp 1681620392
transform 1 0 1076 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5158
timestamp 1681620392
transform 1 0 1164 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5159
timestamp 1681620392
transform 1 0 1188 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5226
timestamp 1681620392
transform 1 0 1076 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5227
timestamp 1681620392
transform 1 0 1116 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5228
timestamp 1681620392
transform 1 0 1180 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4535
timestamp 1681620392
transform 1 0 1060 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4467
timestamp 1681620392
transform 1 0 1220 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4468
timestamp 1681620392
transform 1 0 1276 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_5160
timestamp 1681620392
transform 1 0 1204 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4488
timestamp 1681620392
transform 1 0 1212 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_5161
timestamp 1681620392
transform 1 0 1220 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4489
timestamp 1681620392
transform 1 0 1236 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_5162
timestamp 1681620392
transform 1 0 1252 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5163
timestamp 1681620392
transform 1 0 1340 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5229
timestamp 1681620392
transform 1 0 1212 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5230
timestamp 1681620392
transform 1 0 1228 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5231
timestamp 1681620392
transform 1 0 1236 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4516
timestamp 1681620392
transform 1 0 1252 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_5232
timestamp 1681620392
transform 1 0 1276 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4517
timestamp 1681620392
transform 1 0 1340 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_5233
timestamp 1681620392
transform 1 0 1348 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5234
timestamp 1681620392
transform 1 0 1356 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4536
timestamp 1681620392
transform 1 0 1236 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4537
timestamp 1681620392
transform 1 0 1348 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4577
timestamp 1681620392
transform 1 0 1340 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4562
timestamp 1681620392
transform 1 0 1356 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_4451
timestamp 1681620392
transform 1 0 1380 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_5125
timestamp 1681620392
transform 1 0 1388 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_5164
timestamp 1681620392
transform 1 0 1380 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4518
timestamp 1681620392
transform 1 0 1380 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_4469
timestamp 1681620392
transform 1 0 1412 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4490
timestamp 1681620392
transform 1 0 1428 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_5235
timestamp 1681620392
transform 1 0 1404 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4519
timestamp 1681620392
transform 1 0 1420 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_4470
timestamp 1681620392
transform 1 0 1460 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4491
timestamp 1681620392
transform 1 0 1452 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_5236
timestamp 1681620392
transform 1 0 1436 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5291
timestamp 1681620392
transform 1 0 1396 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_4538
timestamp 1681620392
transform 1 0 1404 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4563
timestamp 1681620392
transform 1 0 1396 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_4520
timestamp 1681620392
transform 1 0 1452 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_5165
timestamp 1681620392
transform 1 0 1492 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5237
timestamp 1681620392
transform 1 0 1468 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4539
timestamp 1681620392
transform 1 0 1436 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_5292
timestamp 1681620392
transform 1 0 1452 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5293
timestamp 1681620392
transform 1 0 1460 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5313
timestamp 1681620392
transform 1 0 1412 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_4578
timestamp 1681620392
transform 1 0 1380 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4564
timestamp 1681620392
transform 1 0 1420 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_5314
timestamp 1681620392
transform 1 0 1444 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_4579
timestamp 1681620392
transform 1 0 1444 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4540
timestamp 1681620392
transform 1 0 1468 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_5294
timestamp 1681620392
transform 1 0 1484 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5315
timestamp 1681620392
transform 1 0 1468 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_4580
timestamp 1681620392
transform 1 0 1468 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4452
timestamp 1681620392
transform 1 0 1524 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_5166
timestamp 1681620392
transform 1 0 1516 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5238
timestamp 1681620392
transform 1 0 1508 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5239
timestamp 1681620392
transform 1 0 1540 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5240
timestamp 1681620392
transform 1 0 1548 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5295
timestamp 1681620392
transform 1 0 1532 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5296
timestamp 1681620392
transform 1 0 1540 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_4471
timestamp 1681620392
transform 1 0 1564 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_5167
timestamp 1681620392
transform 1 0 1564 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5241
timestamp 1681620392
transform 1 0 1572 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4541
timestamp 1681620392
transform 1 0 1556 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4565
timestamp 1681620392
transform 1 0 1572 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_5126
timestamp 1681620392
transform 1 0 1596 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_5242
timestamp 1681620392
transform 1 0 1596 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5243
timestamp 1681620392
transform 1 0 1604 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4542
timestamp 1681620392
transform 1 0 1596 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4566
timestamp 1681620392
transform 1 0 1596 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_4492
timestamp 1681620392
transform 1 0 1612 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_4521
timestamp 1681620392
transform 1 0 1612 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_5168
timestamp 1681620392
transform 1 0 1636 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4493
timestamp 1681620392
transform 1 0 1644 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_5244
timestamp 1681620392
transform 1 0 1620 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5245
timestamp 1681620392
transform 1 0 1628 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5297
timestamp 1681620392
transform 1 0 1620 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_4543
timestamp 1681620392
transform 1 0 1628 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_5246
timestamp 1681620392
transform 1 0 1652 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5298
timestamp 1681620392
transform 1 0 1636 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5299
timestamp 1681620392
transform 1 0 1668 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5316
timestamp 1681620392
transform 1 0 1660 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_4544
timestamp 1681620392
transform 1 0 1676 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_5247
timestamp 1681620392
transform 1 0 1700 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5169
timestamp 1681620392
transform 1 0 1716 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4433
timestamp 1681620392
transform 1 0 1820 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_4453
timestamp 1681620392
transform 1 0 1788 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_4494
timestamp 1681620392
transform 1 0 1796 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_5170
timestamp 1681620392
transform 1 0 1820 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5248
timestamp 1681620392
transform 1 0 1740 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5249
timestamp 1681620392
transform 1 0 1796 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4472
timestamp 1681620392
transform 1 0 1852 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4473
timestamp 1681620392
transform 1 0 1876 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_5171
timestamp 1681620392
transform 1 0 1852 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4495
timestamp 1681620392
transform 1 0 1860 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_4434
timestamp 1681620392
transform 1 0 1892 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_5172
timestamp 1681620392
transform 1 0 1868 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5173
timestamp 1681620392
transform 1 0 1884 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5250
timestamp 1681620392
transform 1 0 1860 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4567
timestamp 1681620392
transform 1 0 1860 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_4454
timestamp 1681620392
transform 1 0 1908 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_4474
timestamp 1681620392
transform 1 0 1932 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_5174
timestamp 1681620392
transform 1 0 1916 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4496
timestamp 1681620392
transform 1 0 1924 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_5175
timestamp 1681620392
transform 1 0 1932 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5251
timestamp 1681620392
transform 1 0 1900 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5252
timestamp 1681620392
transform 1 0 1908 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5253
timestamp 1681620392
transform 1 0 1924 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4545
timestamp 1681620392
transform 1 0 1908 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4435
timestamp 1681620392
transform 1 0 1948 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_4475
timestamp 1681620392
transform 1 0 1956 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4568
timestamp 1681620392
transform 1 0 1964 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_4476
timestamp 1681620392
transform 1 0 2036 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4477
timestamp 1681620392
transform 1 0 2052 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4478
timestamp 1681620392
transform 1 0 2076 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_5176
timestamp 1681620392
transform 1 0 1988 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4497
timestamp 1681620392
transform 1 0 2020 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_4498
timestamp 1681620392
transform 1 0 2036 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_4499
timestamp 1681620392
transform 1 0 2060 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_4522
timestamp 1681620392
transform 1 0 1988 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_4523
timestamp 1681620392
transform 1 0 2012 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_5254
timestamp 1681620392
transform 1 0 2036 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5255
timestamp 1681620392
transform 1 0 2084 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4436
timestamp 1681620392
transform 1 0 2108 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_4437
timestamp 1681620392
transform 1 0 2124 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_5177
timestamp 1681620392
transform 1 0 2108 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4500
timestamp 1681620392
transform 1 0 2156 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_5256
timestamp 1681620392
transform 1 0 2156 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4479
timestamp 1681620392
transform 1 0 2196 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_5178
timestamp 1681620392
transform 1 0 2204 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5257
timestamp 1681620392
transform 1 0 2196 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5258
timestamp 1681620392
transform 1 0 2204 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4546
timestamp 1681620392
transform 1 0 2204 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4438
timestamp 1681620392
transform 1 0 2252 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_4480
timestamp 1681620392
transform 1 0 2252 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4501
timestamp 1681620392
transform 1 0 2244 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_5179
timestamp 1681620392
transform 1 0 2284 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4547
timestamp 1681620392
transform 1 0 2284 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_5300
timestamp 1681620392
transform 1 0 2292 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_4481
timestamp 1681620392
transform 1 0 2316 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_5180
timestamp 1681620392
transform 1 0 2316 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4439
timestamp 1681620392
transform 1 0 2420 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_4482
timestamp 1681620392
transform 1 0 2412 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_5181
timestamp 1681620392
transform 1 0 2332 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5182
timestamp 1681620392
transform 1 0 2420 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5259
timestamp 1681620392
transform 1 0 2356 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5260
timestamp 1681620392
transform 1 0 2412 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4548
timestamp 1681620392
transform 1 0 2356 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4483
timestamp 1681620392
transform 1 0 2436 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_5183
timestamp 1681620392
transform 1 0 2436 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4524
timestamp 1681620392
transform 1 0 2436 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_5261
timestamp 1681620392
transform 1 0 2444 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5301
timestamp 1681620392
transform 1 0 2436 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_4569
timestamp 1681620392
transform 1 0 2444 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_4525
timestamp 1681620392
transform 1 0 2460 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_5302
timestamp 1681620392
transform 1 0 2460 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5184
timestamp 1681620392
transform 1 0 2484 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4526
timestamp 1681620392
transform 1 0 2492 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_5262
timestamp 1681620392
transform 1 0 2500 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4581
timestamp 1681620392
transform 1 0 2500 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_5185
timestamp 1681620392
transform 1 0 2532 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5186
timestamp 1681620392
transform 1 0 2548 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5187
timestamp 1681620392
transform 1 0 2644 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5263
timestamp 1681620392
transform 1 0 2532 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5264
timestamp 1681620392
transform 1 0 2580 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5265
timestamp 1681620392
transform 1 0 2628 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5266
timestamp 1681620392
transform 1 0 2636 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4549
timestamp 1681620392
transform 1 0 2636 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4582
timestamp 1681620392
transform 1 0 2540 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4583
timestamp 1681620392
transform 1 0 2596 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_5303
timestamp 1681620392
transform 1 0 2652 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_4570
timestamp 1681620392
transform 1 0 2652 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_4440
timestamp 1681620392
transform 1 0 2668 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_5188
timestamp 1681620392
transform 1 0 2668 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4502
timestamp 1681620392
transform 1 0 2676 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_5189
timestamp 1681620392
transform 1 0 2692 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5267
timestamp 1681620392
transform 1 0 2684 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5268
timestamp 1681620392
transform 1 0 2692 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4441
timestamp 1681620392
transform 1 0 2724 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_4455
timestamp 1681620392
transform 1 0 2708 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_4456
timestamp 1681620392
transform 1 0 2756 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_5190
timestamp 1681620392
transform 1 0 2716 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5191
timestamp 1681620392
transform 1 0 2724 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5192
timestamp 1681620392
transform 1 0 2740 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5193
timestamp 1681620392
transform 1 0 2756 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5269
timestamp 1681620392
transform 1 0 2716 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5270
timestamp 1681620392
transform 1 0 2748 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4550
timestamp 1681620392
transform 1 0 2716 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4571
timestamp 1681620392
transform 1 0 2748 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_5194
timestamp 1681620392
transform 1 0 2788 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_4503
timestamp 1681620392
transform 1 0 2812 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_5271
timestamp 1681620392
transform 1 0 2812 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5272
timestamp 1681620392
transform 1 0 2868 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5273
timestamp 1681620392
transform 1 0 2876 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_4551
timestamp 1681620392
transform 1 0 2876 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4572
timestamp 1681620392
transform 1 0 2868 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_4442
timestamp 1681620392
transform 1 0 2900 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_5127
timestamp 1681620392
transform 1 0 2900 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_5195
timestamp 1681620392
transform 1 0 2892 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5196
timestamp 1681620392
transform 1 0 2940 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5274
timestamp 1681620392
transform 1 0 2916 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5304
timestamp 1681620392
transform 1 0 2908 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_4552
timestamp 1681620392
transform 1 0 2916 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_5275
timestamp 1681620392
transform 1 0 2956 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5305
timestamp 1681620392
transform 1 0 2932 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5306
timestamp 1681620392
transform 1 0 2940 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5317
timestamp 1681620392
transform 1 0 2908 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_4443
timestamp 1681620392
transform 1 0 2972 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_5197
timestamp 1681620392
transform 1 0 2972 0 1 335
box -2 -2 2 2
use Project_Top_VIA0  Project_Top_VIA0_54
timestamp 1681620392
transform 1 0 24 0 1 270
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_280
timestamp 1681620392
transform 1 0 72 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_281
timestamp 1681620392
transform 1 0 168 0 -1 370
box -8 -3 104 105
use FILL  FILL_1333
timestamp 1681620392
transform 1 0 264 0 -1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_99
timestamp 1681620392
transform -1 0 296 0 -1 370
box -8 -3 32 105
use INVX2  INVX2_339
timestamp 1681620392
transform 1 0 296 0 -1 370
box -9 -3 26 105
use OAI22X1  OAI22X1_112
timestamp 1681620392
transform -1 0 352 0 -1 370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_282
timestamp 1681620392
transform 1 0 352 0 -1 370
box -8 -3 104 105
use AOI21X1  AOI21X1_39
timestamp 1681620392
transform -1 0 480 0 -1 370
box -7 -3 39 105
use NAND2X1  NAND2X1_295
timestamp 1681620392
transform -1 0 504 0 -1 370
box -8 -3 32 105
use NAND3X1  NAND3X1_106
timestamp 1681620392
transform 1 0 504 0 -1 370
box -8 -3 40 105
use AND2X2  AND2X2_28
timestamp 1681620392
transform 1 0 536 0 -1 370
box -8 -3 40 105
use INVX2  INVX2_340
timestamp 1681620392
transform 1 0 568 0 -1 370
box -9 -3 26 105
use FILL  FILL_1334
timestamp 1681620392
transform 1 0 584 0 -1 370
box -8 -3 16 105
use FILL  FILL_1335
timestamp 1681620392
transform 1 0 592 0 -1 370
box -8 -3 16 105
use FILL  FILL_1336
timestamp 1681620392
transform 1 0 600 0 -1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_107
timestamp 1681620392
transform 1 0 608 0 -1 370
box -8 -3 40 105
use INVX2  INVX2_341
timestamp 1681620392
transform 1 0 640 0 -1 370
box -9 -3 26 105
use NOR2X1  NOR2X1_100
timestamp 1681620392
transform -1 0 680 0 -1 370
box -8 -3 32 105
use INVX2  INVX2_342
timestamp 1681620392
transform 1 0 680 0 -1 370
box -9 -3 26 105
use NAND3X1  NAND3X1_108
timestamp 1681620392
transform 1 0 696 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_109
timestamp 1681620392
transform -1 0 760 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_110
timestamp 1681620392
transform 1 0 760 0 -1 370
box -8 -3 40 105
use FILL  FILL_1337
timestamp 1681620392
transform 1 0 792 0 -1 370
box -8 -3 16 105
use FILL  FILL_1338
timestamp 1681620392
transform 1 0 800 0 -1 370
box -8 -3 16 105
use AND2X2  AND2X2_29
timestamp 1681620392
transform 1 0 808 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_111
timestamp 1681620392
transform 1 0 840 0 -1 370
box -8 -3 40 105
use OAI21X1  OAI21X1_290
timestamp 1681620392
transform 1 0 872 0 -1 370
box -8 -3 34 105
use OAI22X1  OAI22X1_113
timestamp 1681620392
transform -1 0 944 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_114
timestamp 1681620392
transform -1 0 984 0 -1 370
box -8 -3 46 105
use FILL  FILL_1339
timestamp 1681620392
transform 1 0 984 0 -1 370
box -8 -3 16 105
use FILL  FILL_1340
timestamp 1681620392
transform 1 0 992 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_343
timestamp 1681620392
transform -1 0 1016 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_344
timestamp 1681620392
transform -1 0 1032 0 -1 370
box -9 -3 26 105
use OAI21X1  OAI21X1_291
timestamp 1681620392
transform -1 0 1064 0 -1 370
box -8 -3 34 105
use INVX2  INVX2_345
timestamp 1681620392
transform -1 0 1080 0 -1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_283
timestamp 1681620392
transform -1 0 1176 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_346
timestamp 1681620392
transform -1 0 1192 0 -1 370
box -9 -3 26 105
use FILL  FILL_1341
timestamp 1681620392
transform 1 0 1192 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_4589
timestamp 1681620392
transform 1 0 1220 0 1 275
box -3 -3 3 3
use OAI22X1  OAI22X1_115
timestamp 1681620392
transform -1 0 1240 0 -1 370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_284
timestamp 1681620392
transform 1 0 1240 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_347
timestamp 1681620392
transform 1 0 1336 0 -1 370
box -9 -3 26 105
use FILL  FILL_1342
timestamp 1681620392
transform 1 0 1352 0 -1 370
box -8 -3 16 105
use FILL  FILL_1343
timestamp 1681620392
transform 1 0 1360 0 -1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_101
timestamp 1681620392
transform -1 0 1392 0 -1 370
box -8 -3 32 105
use NAND3X1  NAND3X1_112
timestamp 1681620392
transform 1 0 1392 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_113
timestamp 1681620392
transform 1 0 1424 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_115
timestamp 1681620392
transform 1 0 1456 0 -1 370
box -8 -3 40 105
use M3_M2  M3_M2_4590
timestamp 1681620392
transform 1 0 1516 0 1 275
box -3 -3 3 3
use INVX2  INVX2_348
timestamp 1681620392
transform 1 0 1488 0 -1 370
box -9 -3 26 105
use FILL  FILL_1344
timestamp 1681620392
transform 1 0 1504 0 -1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_298
timestamp 1681620392
transform 1 0 1512 0 -1 370
box -8 -3 32 105
use FILL  FILL_1348
timestamp 1681620392
transform 1 0 1536 0 -1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_300
timestamp 1681620392
transform -1 0 1568 0 -1 370
box -8 -3 32 105
use M3_M2  M3_M2_4591
timestamp 1681620392
transform 1 0 1580 0 1 275
box -3 -3 3 3
use AOI21X1  AOI21X1_40
timestamp 1681620392
transform 1 0 1568 0 -1 370
box -7 -3 39 105
use INVX2  INVX2_349
timestamp 1681620392
transform 1 0 1600 0 -1 370
box -9 -3 26 105
use NAND2X1  NAND2X1_301
timestamp 1681620392
transform -1 0 1640 0 -1 370
box -8 -3 32 105
use M3_M2  M3_M2_4592
timestamp 1681620392
transform 1 0 1652 0 1 275
box -3 -3 3 3
use NAND3X1  NAND3X1_116
timestamp 1681620392
transform 1 0 1640 0 -1 370
box -8 -3 40 105
use FILL  FILL_1349
timestamp 1681620392
transform 1 0 1672 0 -1 370
box -8 -3 16 105
use FILL  FILL_1356
timestamp 1681620392
transform 1 0 1680 0 -1 370
box -8 -3 16 105
use FILL  FILL_1357
timestamp 1681620392
transform 1 0 1688 0 -1 370
box -8 -3 16 105
use BUFX2  BUFX2_49
timestamp 1681620392
transform 1 0 1696 0 -1 370
box -5 -3 28 105
use FILL  FILL_1358
timestamp 1681620392
transform 1 0 1720 0 -1 370
box -8 -3 16 105
use FILL  FILL_1359
timestamp 1681620392
transform 1 0 1728 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_286
timestamp 1681620392
transform -1 0 1832 0 -1 370
box -8 -3 104 105
use FILL  FILL_1360
timestamp 1681620392
transform 1 0 1832 0 -1 370
box -8 -3 16 105
use FILL  FILL_1363
timestamp 1681620392
transform 1 0 1840 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_117
timestamp 1681620392
transform -1 0 1888 0 -1 370
box -8 -3 46 105
use FILL  FILL_1364
timestamp 1681620392
transform 1 0 1888 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_119
timestamp 1681620392
transform 1 0 1896 0 -1 370
box -8 -3 46 105
use FILL  FILL_1372
timestamp 1681620392
transform 1 0 1936 0 -1 370
box -8 -3 16 105
use FILL  FILL_1373
timestamp 1681620392
transform 1 0 1944 0 -1 370
box -8 -3 16 105
use FILL  FILL_1374
timestamp 1681620392
transform 1 0 1952 0 -1 370
box -8 -3 16 105
use FILL  FILL_1375
timestamp 1681620392
transform 1 0 1960 0 -1 370
box -8 -3 16 105
use FILL  FILL_1376
timestamp 1681620392
transform 1 0 1968 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_289
timestamp 1681620392
transform 1 0 1976 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_351
timestamp 1681620392
transform 1 0 2072 0 -1 370
box -9 -3 26 105
use FILL  FILL_1377
timestamp 1681620392
transform 1 0 2088 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_290
timestamp 1681620392
transform 1 0 2096 0 -1 370
box -8 -3 104 105
use FILL  FILL_1378
timestamp 1681620392
transform 1 0 2192 0 -1 370
box -8 -3 16 105
use FILL  FILL_1379
timestamp 1681620392
transform 1 0 2200 0 -1 370
box -8 -3 16 105
use FILL  FILL_1380
timestamp 1681620392
transform 1 0 2208 0 -1 370
box -8 -3 16 105
use FILL  FILL_1381
timestamp 1681620392
transform 1 0 2216 0 -1 370
box -8 -3 16 105
use FILL  FILL_1382
timestamp 1681620392
transform 1 0 2224 0 -1 370
box -8 -3 16 105
use FILL  FILL_1383
timestamp 1681620392
transform 1 0 2232 0 -1 370
box -8 -3 16 105
use FILL  FILL_1384
timestamp 1681620392
transform 1 0 2240 0 -1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_297
timestamp 1681620392
transform 1 0 2248 0 -1 370
box -8 -3 34 105
use FILL  FILL_1385
timestamp 1681620392
transform 1 0 2280 0 -1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_305
timestamp 1681620392
transform -1 0 2312 0 -1 370
box -8 -3 32 105
use FILL  FILL_1386
timestamp 1681620392
transform 1 0 2312 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_292
timestamp 1681620392
transform 1 0 2320 0 -1 370
box -8 -3 104 105
use NAND2X1  NAND2X1_307
timestamp 1681620392
transform 1 0 2416 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_308
timestamp 1681620392
transform 1 0 2440 0 -1 370
box -8 -3 32 105
use FILL  FILL_1396
timestamp 1681620392
transform 1 0 2464 0 -1 370
box -8 -3 16 105
use FILL  FILL_1397
timestamp 1681620392
transform 1 0 2472 0 -1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_299
timestamp 1681620392
transform -1 0 2512 0 -1 370
box -8 -3 34 105
use FILL  FILL_1398
timestamp 1681620392
transform 1 0 2512 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_353
timestamp 1681620392
transform -1 0 2536 0 -1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_294
timestamp 1681620392
transform 1 0 2536 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_354
timestamp 1681620392
transform -1 0 2648 0 -1 370
box -9 -3 26 105
use FILL  FILL_1399
timestamp 1681620392
transform 1 0 2648 0 -1 370
box -8 -3 16 105
use FILL  FILL_1404
timestamp 1681620392
transform 1 0 2656 0 -1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_300
timestamp 1681620392
transform -1 0 2696 0 -1 370
box -8 -3 34 105
use FILL  FILL_1405
timestamp 1681620392
transform 1 0 2696 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_355
timestamp 1681620392
transform -1 0 2720 0 -1 370
box -9 -3 26 105
use OAI22X1  OAI22X1_121
timestamp 1681620392
transform 1 0 2720 0 -1 370
box -8 -3 46 105
use FILL  FILL_1406
timestamp 1681620392
transform 1 0 2760 0 -1 370
box -8 -3 16 105
use FILL  FILL_1408
timestamp 1681620392
transform 1 0 2768 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_295
timestamp 1681620392
transform 1 0 2776 0 -1 370
box -8 -3 104 105
use FILL  FILL_1419
timestamp 1681620392
transform 1 0 2872 0 -1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_102
timestamp 1681620392
transform -1 0 2904 0 -1 370
box -8 -3 32 105
use NAND3X1  NAND3X1_117
timestamp 1681620392
transform 1 0 2904 0 -1 370
box -8 -3 40 105
use OAI21X1  OAI21X1_303
timestamp 1681620392
transform -1 0 2968 0 -1 370
box -8 -3 34 105
use FILL  FILL_1420
timestamp 1681620392
transform 1 0 2968 0 -1 370
box -8 -3 16 105
use FILL  FILL_1422
timestamp 1681620392
transform 1 0 2976 0 -1 370
box -8 -3 16 105
use FILL  FILL_1424
timestamp 1681620392
transform 1 0 2984 0 -1 370
box -8 -3 16 105
use FILL  FILL_1426
timestamp 1681620392
transform 1 0 2992 0 -1 370
box -8 -3 16 105
use FILL  FILL_1428
timestamp 1681620392
transform 1 0 3000 0 -1 370
box -8 -3 16 105
use FILL  FILL_1430
timestamp 1681620392
transform 1 0 3008 0 -1 370
box -8 -3 16 105
use Project_Top_VIA0  Project_Top_VIA0_55
timestamp 1681620392
transform 1 0 3067 0 1 270
box -10 -3 10 3
use M3_M2  M3_M2_4613
timestamp 1681620392
transform 1 0 204 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_4614
timestamp 1681620392
transform 1 0 236 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_4630
timestamp 1681620392
transform 1 0 164 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5363
timestamp 1681620392
transform 1 0 132 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5364
timestamp 1681620392
transform 1 0 164 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5365
timestamp 1681620392
transform 1 0 180 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5366
timestamp 1681620392
transform 1 0 204 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4667
timestamp 1681620392
transform 1 0 212 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_4631
timestamp 1681620392
transform 1 0 260 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5367
timestamp 1681620392
transform 1 0 220 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5368
timestamp 1681620392
transform 1 0 236 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5369
timestamp 1681620392
transform 1 0 244 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5450
timestamp 1681620392
transform 1 0 84 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5451
timestamp 1681620392
transform 1 0 172 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4696
timestamp 1681620392
transform 1 0 132 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4690
timestamp 1681620392
transform 1 0 180 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_5452
timestamp 1681620392
transform 1 0 188 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5453
timestamp 1681620392
transform 1 0 204 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5454
timestamp 1681620392
transform 1 0 212 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5455
timestamp 1681620392
transform 1 0 228 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5456
timestamp 1681620392
transform 1 0 244 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5457
timestamp 1681620392
transform 1 0 260 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4726
timestamp 1681620392
transform 1 0 172 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_4697
timestamp 1681620392
transform 1 0 228 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4727
timestamp 1681620392
transform 1 0 212 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_5535
timestamp 1681620392
transform 1 0 268 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_4597
timestamp 1681620392
transform 1 0 300 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_4601
timestamp 1681620392
transform 1 0 292 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_4632
timestamp 1681620392
transform 1 0 284 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5370
timestamp 1681620392
transform 1 0 284 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4615
timestamp 1681620392
transform 1 0 308 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_5371
timestamp 1681620392
transform 1 0 308 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4668
timestamp 1681620392
transform 1 0 316 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_5458
timestamp 1681620392
transform 1 0 292 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5459
timestamp 1681620392
transform 1 0 300 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5536
timestamp 1681620392
transform 1 0 284 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_5460
timestamp 1681620392
transform 1 0 316 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4616
timestamp 1681620392
transform 1 0 348 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_4633
timestamp 1681620392
transform 1 0 332 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5372
timestamp 1681620392
transform 1 0 332 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5373
timestamp 1681620392
transform 1 0 348 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5461
timestamp 1681620392
transform 1 0 340 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5462
timestamp 1681620392
transform 1 0 388 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4634
timestamp 1681620392
transform 1 0 404 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5374
timestamp 1681620392
transform 1 0 412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5537
timestamp 1681620392
transform 1 0 404 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_4635
timestamp 1681620392
transform 1 0 436 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5375
timestamp 1681620392
transform 1 0 428 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5376
timestamp 1681620392
transform 1 0 436 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5463
timestamp 1681620392
transform 1 0 420 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5377
timestamp 1681620392
transform 1 0 468 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5464
timestamp 1681620392
transform 1 0 444 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5465
timestamp 1681620392
transform 1 0 460 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4698
timestamp 1681620392
transform 1 0 420 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_5466
timestamp 1681620392
transform 1 0 476 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4699
timestamp 1681620392
transform 1 0 476 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4602
timestamp 1681620392
transform 1 0 516 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_5318
timestamp 1681620392
transform 1 0 524 0 1 235
box -2 -2 2 2
use M3_M2  M3_M2_4636
timestamp 1681620392
transform 1 0 508 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5327
timestamp 1681620392
transform 1 0 516 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5328
timestamp 1681620392
transform 1 0 532 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5378
timestamp 1681620392
transform 1 0 508 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4637
timestamp 1681620392
transform 1 0 540 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5329
timestamp 1681620392
transform 1 0 556 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_4638
timestamp 1681620392
transform 1 0 564 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5379
timestamp 1681620392
transform 1 0 532 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4669
timestamp 1681620392
transform 1 0 556 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_5330
timestamp 1681620392
transform 1 0 604 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5331
timestamp 1681620392
transform 1 0 612 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5380
timestamp 1681620392
transform 1 0 564 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5381
timestamp 1681620392
transform 1 0 588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5382
timestamp 1681620392
transform 1 0 596 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5467
timestamp 1681620392
transform 1 0 556 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4700
timestamp 1681620392
transform 1 0 540 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_5468
timestamp 1681620392
transform 1 0 588 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4598
timestamp 1681620392
transform 1 0 628 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_5383
timestamp 1681620392
transform 1 0 620 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5384
timestamp 1681620392
transform 1 0 628 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5469
timestamp 1681620392
transform 1 0 636 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5332
timestamp 1681620392
transform 1 0 652 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_4639
timestamp 1681620392
transform 1 0 660 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5385
timestamp 1681620392
transform 1 0 660 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5470
timestamp 1681620392
transform 1 0 652 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4593
timestamp 1681620392
transform 1 0 676 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_4603
timestamp 1681620392
transform 1 0 676 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_4594
timestamp 1681620392
transform 1 0 716 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_4604
timestamp 1681620392
transform 1 0 708 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_5319
timestamp 1681620392
transform 1 0 700 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_5333
timestamp 1681620392
transform 1 0 676 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5334
timestamp 1681620392
transform 1 0 684 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5335
timestamp 1681620392
transform 1 0 692 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5336
timestamp 1681620392
transform 1 0 708 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5337
timestamp 1681620392
transform 1 0 716 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5386
timestamp 1681620392
transform 1 0 676 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5471
timestamp 1681620392
transform 1 0 692 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4701
timestamp 1681620392
transform 1 0 692 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4595
timestamp 1681620392
transform 1 0 756 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_4640
timestamp 1681620392
transform 1 0 764 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5387
timestamp 1681620392
transform 1 0 724 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5388
timestamp 1681620392
transform 1 0 732 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5389
timestamp 1681620392
transform 1 0 748 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5472
timestamp 1681620392
transform 1 0 732 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4702
timestamp 1681620392
transform 1 0 724 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_5390
timestamp 1681620392
transform 1 0 788 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5391
timestamp 1681620392
transform 1 0 796 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5473
timestamp 1681620392
transform 1 0 764 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5474
timestamp 1681620392
transform 1 0 772 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5538
timestamp 1681620392
transform 1 0 788 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_4596
timestamp 1681620392
transform 1 0 820 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_5320
timestamp 1681620392
transform 1 0 828 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_5338
timestamp 1681620392
transform 1 0 812 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_4641
timestamp 1681620392
transform 1 0 828 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5339
timestamp 1681620392
transform 1 0 836 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5340
timestamp 1681620392
transform 1 0 844 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5392
timestamp 1681620392
transform 1 0 820 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5475
timestamp 1681620392
transform 1 0 804 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4703
timestamp 1681620392
transform 1 0 804 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4670
timestamp 1681620392
transform 1 0 844 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_4642
timestamp 1681620392
transform 1 0 868 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5321
timestamp 1681620392
transform 1 0 916 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_5341
timestamp 1681620392
transform 1 0 892 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5342
timestamp 1681620392
transform 1 0 900 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_4643
timestamp 1681620392
transform 1 0 908 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5393
timestamp 1681620392
transform 1 0 876 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5394
timestamp 1681620392
transform 1 0 884 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5476
timestamp 1681620392
transform 1 0 860 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5477
timestamp 1681620392
transform 1 0 868 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4671
timestamp 1681620392
transform 1 0 892 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_5395
timestamp 1681620392
transform 1 0 908 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4672
timestamp 1681620392
transform 1 0 916 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_4605
timestamp 1681620392
transform 1 0 948 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_5478
timestamp 1681620392
transform 1 0 948 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5343
timestamp 1681620392
transform 1 0 956 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5396
timestamp 1681620392
transform 1 0 972 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5397
timestamp 1681620392
transform 1 0 996 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5398
timestamp 1681620392
transform 1 0 1036 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5399
timestamp 1681620392
transform 1 0 1092 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5479
timestamp 1681620392
transform 1 0 980 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5480
timestamp 1681620392
transform 1 0 996 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5481
timestamp 1681620392
transform 1 0 1012 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4704
timestamp 1681620392
transform 1 0 980 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4705
timestamp 1681620392
transform 1 0 1036 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4728
timestamp 1681620392
transform 1 0 1012 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_4644
timestamp 1681620392
transform 1 0 1108 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5400
timestamp 1681620392
transform 1 0 1108 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4729
timestamp 1681620392
transform 1 0 1108 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_4617
timestamp 1681620392
transform 1 0 1132 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_4645
timestamp 1681620392
transform 1 0 1148 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5401
timestamp 1681620392
transform 1 0 1116 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5402
timestamp 1681620392
transform 1 0 1132 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5403
timestamp 1681620392
transform 1 0 1148 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5482
timestamp 1681620392
transform 1 0 1124 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5483
timestamp 1681620392
transform 1 0 1140 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5484
timestamp 1681620392
transform 1 0 1156 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4706
timestamp 1681620392
transform 1 0 1124 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4646
timestamp 1681620392
transform 1 0 1196 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5404
timestamp 1681620392
transform 1 0 1180 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5405
timestamp 1681620392
transform 1 0 1196 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5485
timestamp 1681620392
transform 1 0 1172 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4691
timestamp 1681620392
transform 1 0 1180 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_4647
timestamp 1681620392
transform 1 0 1228 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_4648
timestamp 1681620392
transform 1 0 1244 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_4649
timestamp 1681620392
transform 1 0 1356 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5406
timestamp 1681620392
transform 1 0 1220 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5407
timestamp 1681620392
transform 1 0 1236 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5408
timestamp 1681620392
transform 1 0 1244 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5409
timestamp 1681620392
transform 1 0 1284 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5410
timestamp 1681620392
transform 1 0 1348 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5411
timestamp 1681620392
transform 1 0 1356 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5486
timestamp 1681620392
transform 1 0 1188 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5487
timestamp 1681620392
transform 1 0 1204 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5488
timestamp 1681620392
transform 1 0 1212 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5489
timestamp 1681620392
transform 1 0 1228 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4707
timestamp 1681620392
transform 1 0 1172 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4730
timestamp 1681620392
transform 1 0 1164 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_4708
timestamp 1681620392
transform 1 0 1212 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4709
timestamp 1681620392
transform 1 0 1228 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_5490
timestamp 1681620392
transform 1 0 1260 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5491
timestamp 1681620392
transform 1 0 1348 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4710
timestamp 1681620392
transform 1 0 1284 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4618
timestamp 1681620392
transform 1 0 1380 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_5412
timestamp 1681620392
transform 1 0 1372 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5492
timestamp 1681620392
transform 1 0 1364 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4711
timestamp 1681620392
transform 1 0 1364 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4731
timestamp 1681620392
transform 1 0 1372 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_4599
timestamp 1681620392
transform 1 0 1428 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_5322
timestamp 1681620392
transform 1 0 1420 0 1 235
box -2 -2 2 2
use M3_M2  M3_M2_4600
timestamp 1681620392
transform 1 0 1460 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_5323
timestamp 1681620392
transform 1 0 1452 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_5344
timestamp 1681620392
transform 1 0 1396 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5345
timestamp 1681620392
transform 1 0 1404 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5346
timestamp 1681620392
transform 1 0 1428 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_4673
timestamp 1681620392
transform 1 0 1396 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_4650
timestamp 1681620392
transform 1 0 1444 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_4606
timestamp 1681620392
transform 1 0 1476 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_5347
timestamp 1681620392
transform 1 0 1460 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_4674
timestamp 1681620392
transform 1 0 1428 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_5413
timestamp 1681620392
transform 1 0 1444 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5493
timestamp 1681620392
transform 1 0 1396 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5494
timestamp 1681620392
transform 1 0 1412 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4712
timestamp 1681620392
transform 1 0 1412 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_5495
timestamp 1681620392
transform 1 0 1468 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5348
timestamp 1681620392
transform 1 0 1484 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_4607
timestamp 1681620392
transform 1 0 1500 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_5414
timestamp 1681620392
transform 1 0 1492 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4608
timestamp 1681620392
transform 1 0 1540 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_4619
timestamp 1681620392
transform 1 0 1532 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_5324
timestamp 1681620392
transform 1 0 1540 0 1 235
box -2 -2 2 2
use M3_M2  M3_M2_4620
timestamp 1681620392
transform 1 0 1548 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_4651
timestamp 1681620392
transform 1 0 1508 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_4652
timestamp 1681620392
transform 1 0 1524 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5349
timestamp 1681620392
transform 1 0 1532 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5350
timestamp 1681620392
transform 1 0 1548 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5415
timestamp 1681620392
transform 1 0 1508 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5416
timestamp 1681620392
transform 1 0 1524 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5417
timestamp 1681620392
transform 1 0 1548 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5496
timestamp 1681620392
transform 1 0 1500 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4713
timestamp 1681620392
transform 1 0 1492 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4732
timestamp 1681620392
transform 1 0 1484 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_4621
timestamp 1681620392
transform 1 0 1588 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_5325
timestamp 1681620392
transform 1 0 1596 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_5326
timestamp 1681620392
transform 1 0 1604 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_5351
timestamp 1681620392
transform 1 0 1588 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_4675
timestamp 1681620392
transform 1 0 1572 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_5418
timestamp 1681620392
transform 1 0 1580 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4676
timestamp 1681620392
transform 1 0 1588 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_5352
timestamp 1681620392
transform 1 0 1612 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5419
timestamp 1681620392
transform 1 0 1596 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5497
timestamp 1681620392
transform 1 0 1564 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5539
timestamp 1681620392
transform 1 0 1564 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_4677
timestamp 1681620392
transform 1 0 1612 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_4733
timestamp 1681620392
transform 1 0 1604 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_5353
timestamp 1681620392
transform 1 0 1644 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_4678
timestamp 1681620392
transform 1 0 1636 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_5420
timestamp 1681620392
transform 1 0 1652 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5421
timestamp 1681620392
transform 1 0 1668 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5498
timestamp 1681620392
transform 1 0 1636 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5499
timestamp 1681620392
transform 1 0 1644 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4714
timestamp 1681620392
transform 1 0 1644 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4653
timestamp 1681620392
transform 1 0 1884 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_4679
timestamp 1681620392
transform 1 0 1836 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_5422
timestamp 1681620392
transform 1 0 1844 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5423
timestamp 1681620392
transform 1 0 1884 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5500
timestamp 1681620392
transform 1 0 1796 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5501
timestamp 1681620392
transform 1 0 1884 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4609
timestamp 1681620392
transform 1 0 1892 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_4654
timestamp 1681620392
transform 1 0 1900 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5424
timestamp 1681620392
transform 1 0 1892 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5425
timestamp 1681620392
transform 1 0 1900 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5426
timestamp 1681620392
transform 1 0 1908 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4680
timestamp 1681620392
transform 1 0 1916 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_5427
timestamp 1681620392
transform 1 0 1924 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5428
timestamp 1681620392
transform 1 0 1940 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4655
timestamp 1681620392
transform 1 0 1996 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5429
timestamp 1681620392
transform 1 0 1964 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4681
timestamp 1681620392
transform 1 0 1988 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_5430
timestamp 1681620392
transform 1 0 1996 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5502
timestamp 1681620392
transform 1 0 1916 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5503
timestamp 1681620392
transform 1 0 1932 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5504
timestamp 1681620392
transform 1 0 1948 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5505
timestamp 1681620392
transform 1 0 1956 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5506
timestamp 1681620392
transform 1 0 1972 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4715
timestamp 1681620392
transform 1 0 1916 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4692
timestamp 1681620392
transform 1 0 1980 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_5507
timestamp 1681620392
transform 1 0 1988 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4716
timestamp 1681620392
transform 1 0 1956 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4734
timestamp 1681620392
transform 1 0 1948 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_4735
timestamp 1681620392
transform 1 0 1988 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_4622
timestamp 1681620392
transform 1 0 2084 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_5431
timestamp 1681620392
transform 1 0 2036 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4682
timestamp 1681620392
transform 1 0 2052 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_5508
timestamp 1681620392
transform 1 0 2012 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4693
timestamp 1681620392
transform 1 0 2036 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_4736
timestamp 1681620392
transform 1 0 2012 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_4737
timestamp 1681620392
transform 1 0 2084 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_4656
timestamp 1681620392
transform 1 0 2108 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5432
timestamp 1681620392
transform 1 0 2108 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5509
timestamp 1681620392
transform 1 0 2124 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4717
timestamp 1681620392
transform 1 0 2124 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4623
timestamp 1681620392
transform 1 0 2172 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_5354
timestamp 1681620392
transform 1 0 2156 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_4657
timestamp 1681620392
transform 1 0 2164 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5510
timestamp 1681620392
transform 1 0 2148 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5433
timestamp 1681620392
transform 1 0 2172 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5511
timestamp 1681620392
transform 1 0 2172 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5512
timestamp 1681620392
transform 1 0 2180 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4718
timestamp 1681620392
transform 1 0 2180 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4610
timestamp 1681620392
transform 1 0 2252 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_4624
timestamp 1681620392
transform 1 0 2236 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_4658
timestamp 1681620392
transform 1 0 2228 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5355
timestamp 1681620392
transform 1 0 2236 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5513
timestamp 1681620392
transform 1 0 2228 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5434
timestamp 1681620392
transform 1 0 2252 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4625
timestamp 1681620392
transform 1 0 2284 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_5514
timestamp 1681620392
transform 1 0 2276 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4683
timestamp 1681620392
transform 1 0 2292 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_5515
timestamp 1681620392
transform 1 0 2292 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4626
timestamp 1681620392
transform 1 0 2316 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_4627
timestamp 1681620392
transform 1 0 2340 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_5356
timestamp 1681620392
transform 1 0 2316 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5357
timestamp 1681620392
transform 1 0 2324 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_4659
timestamp 1681620392
transform 1 0 2332 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5358
timestamp 1681620392
transform 1 0 2348 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_4684
timestamp 1681620392
transform 1 0 2324 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_5435
timestamp 1681620392
transform 1 0 2332 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5436
timestamp 1681620392
transform 1 0 2340 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4685
timestamp 1681620392
transform 1 0 2348 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_5516
timestamp 1681620392
transform 1 0 2324 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5517
timestamp 1681620392
transform 1 0 2348 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4719
timestamp 1681620392
transform 1 0 2324 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4660
timestamp 1681620392
transform 1 0 2380 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5437
timestamp 1681620392
transform 1 0 2404 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5518
timestamp 1681620392
transform 1 0 2364 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5519
timestamp 1681620392
transform 1 0 2380 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4720
timestamp 1681620392
transform 1 0 2404 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4738
timestamp 1681620392
transform 1 0 2364 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_5520
timestamp 1681620392
transform 1 0 2468 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4739
timestamp 1681620392
transform 1 0 2468 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_4611
timestamp 1681620392
transform 1 0 2508 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_4628
timestamp 1681620392
transform 1 0 2500 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_4629
timestamp 1681620392
transform 1 0 2524 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_5359
timestamp 1681620392
transform 1 0 2492 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5360
timestamp 1681620392
transform 1 0 2516 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5361
timestamp 1681620392
transform 1 0 2524 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_4661
timestamp 1681620392
transform 1 0 2532 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_4686
timestamp 1681620392
transform 1 0 2492 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_5438
timestamp 1681620392
transform 1 0 2500 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5439
timestamp 1681620392
transform 1 0 2508 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4687
timestamp 1681620392
transform 1 0 2516 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_5440
timestamp 1681620392
transform 1 0 2540 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5521
timestamp 1681620392
transform 1 0 2492 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5522
timestamp 1681620392
transform 1 0 2524 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4721
timestamp 1681620392
transform 1 0 2524 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4688
timestamp 1681620392
transform 1 0 2548 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_5441
timestamp 1681620392
transform 1 0 2588 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4689
timestamp 1681620392
transform 1 0 2636 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_4612
timestamp 1681620392
transform 1 0 2652 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_5362
timestamp 1681620392
transform 1 0 2652 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5442
timestamp 1681620392
transform 1 0 2644 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5523
timestamp 1681620392
transform 1 0 2548 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5524
timestamp 1681620392
transform 1 0 2564 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4722
timestamp 1681620392
transform 1 0 2588 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4662
timestamp 1681620392
transform 1 0 2700 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5443
timestamp 1681620392
transform 1 0 2692 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5444
timestamp 1681620392
transform 1 0 2700 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5525
timestamp 1681620392
transform 1 0 2676 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4694
timestamp 1681620392
transform 1 0 2684 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_5445
timestamp 1681620392
transform 1 0 2740 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4663
timestamp 1681620392
transform 1 0 2764 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_4664
timestamp 1681620392
transform 1 0 2788 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5446
timestamp 1681620392
transform 1 0 2788 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5526
timestamp 1681620392
transform 1 0 2708 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5527
timestamp 1681620392
transform 1 0 2716 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5528
timestamp 1681620392
transform 1 0 2732 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5529
timestamp 1681620392
transform 1 0 2748 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5530
timestamp 1681620392
transform 1 0 2764 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_4723
timestamp 1681620392
transform 1 0 2708 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4695
timestamp 1681620392
transform 1 0 2788 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_4724
timestamp 1681620392
transform 1 0 2828 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_5447
timestamp 1681620392
transform 1 0 2860 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5448
timestamp 1681620392
transform 1 0 2868 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4725
timestamp 1681620392
transform 1 0 2860 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4665
timestamp 1681620392
transform 1 0 2892 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_4666
timestamp 1681620392
transform 1 0 2924 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_5531
timestamp 1681620392
transform 1 0 2892 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5532
timestamp 1681620392
transform 1 0 2900 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5540
timestamp 1681620392
transform 1 0 2892 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_5449
timestamp 1681620392
transform 1 0 2924 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_4740
timestamp 1681620392
transform 1 0 2892 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_4741
timestamp 1681620392
transform 1 0 2908 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_5533
timestamp 1681620392
transform 1 0 2940 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5534
timestamp 1681620392
transform 1 0 2972 0 1 205
box -2 -2 2 2
use Project_Top_VIA0  Project_Top_VIA0_56
timestamp 1681620392
transform 1 0 48 0 1 170
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_296
timestamp 1681620392
transform 1 0 72 0 1 170
box -8 -3 104 105
use M3_M2  M3_M2_4742
timestamp 1681620392
transform 1 0 204 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_122
timestamp 1681620392
transform -1 0 208 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_123
timestamp 1681620392
transform -1 0 248 0 1 170
box -8 -3 46 105
use M3_M2  M3_M2_4743
timestamp 1681620392
transform 1 0 268 0 1 175
box -3 -3 3 3
use INVX2  INVX2_358
timestamp 1681620392
transform -1 0 264 0 1 170
box -9 -3 26 105
use NOR2X1  NOR2X1_103
timestamp 1681620392
transform 1 0 264 0 1 170
box -8 -3 32 105
use M3_M2  M3_M2_4744
timestamp 1681620392
transform 1 0 300 0 1 175
box -3 -3 3 3
use NOR2X1  NOR2X1_104
timestamp 1681620392
transform 1 0 288 0 1 170
box -8 -3 32 105
use FILL  FILL_1431
timestamp 1681620392
transform 1 0 312 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_4745
timestamp 1681620392
transform 1 0 364 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_124
timestamp 1681620392
transform -1 0 360 0 1 170
box -8 -3 46 105
use INVX2  INVX2_359
timestamp 1681620392
transform -1 0 376 0 1 170
box -9 -3 26 105
use FILL  FILL_1432
timestamp 1681620392
transform 1 0 376 0 1 170
box -8 -3 16 105
use FILL  FILL_1433
timestamp 1681620392
transform 1 0 384 0 1 170
box -8 -3 16 105
use FILL  FILL_1434
timestamp 1681620392
transform 1 0 392 0 1 170
box -8 -3 16 105
use FILL  FILL_1444
timestamp 1681620392
transform 1 0 400 0 1 170
box -8 -3 16 105
use NOR2X1  NOR2X1_107
timestamp 1681620392
transform 1 0 408 0 1 170
box -8 -3 32 105
use INVX2  INVX2_361
timestamp 1681620392
transform -1 0 448 0 1 170
box -9 -3 26 105
use M3_M2  M3_M2_4746
timestamp 1681620392
transform 1 0 476 0 1 175
box -3 -3 3 3
use NOR2X1  NOR2X1_108
timestamp 1681620392
transform 1 0 448 0 1 170
box -8 -3 32 105
use FILL  FILL_1448
timestamp 1681620392
transform 1 0 472 0 1 170
box -8 -3 16 105
use FILL  FILL_1450
timestamp 1681620392
transform 1 0 480 0 1 170
box -8 -3 16 105
use FILL  FILL_1452
timestamp 1681620392
transform 1 0 488 0 1 170
box -8 -3 16 105
use NAND2X1  NAND2X1_310
timestamp 1681620392
transform 1 0 496 0 1 170
box -8 -3 32 105
use NAND3X1  NAND3X1_118
timestamp 1681620392
transform 1 0 520 0 1 170
box -8 -3 40 105
use M3_M2  M3_M2_4747
timestamp 1681620392
transform 1 0 588 0 1 175
box -3 -3 3 3
use AND2X2  AND2X2_30
timestamp 1681620392
transform 1 0 552 0 1 170
box -8 -3 40 105
use M3_M2  M3_M2_4748
timestamp 1681620392
transform 1 0 612 0 1 175
box -3 -3 3 3
use NAND2X1  NAND2X1_311
timestamp 1681620392
transform 1 0 584 0 1 170
box -8 -3 32 105
use M3_M2  M3_M2_4749
timestamp 1681620392
transform 1 0 628 0 1 175
box -3 -3 3 3
use NAND2X1  NAND2X1_312
timestamp 1681620392
transform -1 0 632 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_313
timestamp 1681620392
transform 1 0 632 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_314
timestamp 1681620392
transform 1 0 656 0 1 170
box -8 -3 32 105
use NAND3X1  NAND3X1_119
timestamp 1681620392
transform 1 0 680 0 1 170
box -8 -3 40 105
use NAND2X1  NAND2X1_315
timestamp 1681620392
transform -1 0 736 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_316
timestamp 1681620392
transform 1 0 736 0 1 170
box -8 -3 32 105
use M3_M2  M3_M2_4750
timestamp 1681620392
transform 1 0 772 0 1 175
box -3 -3 3 3
use AOI21X1  AOI21X1_41
timestamp 1681620392
transform 1 0 760 0 1 170
box -7 -3 39 105
use INVX2  INVX2_362
timestamp 1681620392
transform -1 0 808 0 1 170
box -9 -3 26 105
use NAND3X1  NAND3X1_120
timestamp 1681620392
transform 1 0 808 0 1 170
box -8 -3 40 105
use NAND2X1  NAND2X1_317
timestamp 1681620392
transform -1 0 864 0 1 170
box -8 -3 32 105
use FILL  FILL_1454
timestamp 1681620392
transform 1 0 864 0 1 170
box -8 -3 16 105
use NAND2X1  NAND2X1_318
timestamp 1681620392
transform 1 0 872 0 1 170
box -8 -3 32 105
use NAND3X1  NAND3X1_121
timestamp 1681620392
transform 1 0 896 0 1 170
box -8 -3 40 105
use FILL  FILL_1455
timestamp 1681620392
transform 1 0 928 0 1 170
box -8 -3 16 105
use FILL  FILL_1456
timestamp 1681620392
transform 1 0 936 0 1 170
box -8 -3 16 105
use FILL  FILL_1457
timestamp 1681620392
transform 1 0 944 0 1 170
box -8 -3 16 105
use FILL  FILL_1458
timestamp 1681620392
transform 1 0 952 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_125
timestamp 1681620392
transform -1 0 1000 0 1 170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_299
timestamp 1681620392
transform 1 0 1000 0 1 170
box -8 -3 104 105
use FILL  FILL_1459
timestamp 1681620392
transform 1 0 1096 0 1 170
box -8 -3 16 105
use INVX2  INVX2_363
timestamp 1681620392
transform 1 0 1104 0 1 170
box -9 -3 26 105
use OAI22X1  OAI22X1_126
timestamp 1681620392
transform -1 0 1160 0 1 170
box -8 -3 46 105
use FILL  FILL_1460
timestamp 1681620392
transform 1 0 1160 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_4751
timestamp 1681620392
transform 1 0 1204 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_127
timestamp 1681620392
transform -1 0 1208 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_128
timestamp 1681620392
transform -1 0 1248 0 1 170
box -8 -3 46 105
use M3_M2  M3_M2_4752
timestamp 1681620392
transform 1 0 1340 0 1 175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_300
timestamp 1681620392
transform 1 0 1248 0 1 170
box -8 -3 104 105
use INVX2  INVX2_364
timestamp 1681620392
transform 1 0 1344 0 1 170
box -9 -3 26 105
use FILL  FILL_1461
timestamp 1681620392
transform 1 0 1360 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_304
timestamp 1681620392
transform 1 0 1368 0 1 170
box -8 -3 34 105
use NAND3X1  NAND3X1_122
timestamp 1681620392
transform 1 0 1400 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_123
timestamp 1681620392
transform 1 0 1432 0 1 170
box -8 -3 40 105
use NAND2X1  NAND2X1_319
timestamp 1681620392
transform 1 0 1464 0 1 170
box -8 -3 32 105
use FILL  FILL_1484
timestamp 1681620392
transform 1 0 1488 0 1 170
box -8 -3 16 105
use AND2X2  AND2X2_32
timestamp 1681620392
transform 1 0 1496 0 1 170
box -8 -3 40 105
use M3_M2  M3_M2_4753
timestamp 1681620392
transform 1 0 1548 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_4754
timestamp 1681620392
transform 1 0 1564 0 1 175
box -3 -3 3 3
use NAND3X1  NAND3X1_126
timestamp 1681620392
transform -1 0 1560 0 1 170
box -8 -3 40 105
use NOR2X1  NOR2X1_114
timestamp 1681620392
transform 1 0 1560 0 1 170
box -8 -3 32 105
use M3_M2  M3_M2_4755
timestamp 1681620392
transform 1 0 1596 0 1 175
box -3 -3 3 3
use NAND3X1  NAND3X1_127
timestamp 1681620392
transform 1 0 1584 0 1 170
box -8 -3 40 105
use INVX2  INVX2_372
timestamp 1681620392
transform -1 0 1632 0 1 170
box -9 -3 26 105
use FILL  FILL_1486
timestamp 1681620392
transform 1 0 1632 0 1 170
box -8 -3 16 105
use AND2X2  AND2X2_33
timestamp 1681620392
transform 1 0 1640 0 1 170
box -8 -3 40 105
use FILL  FILL_1494
timestamp 1681620392
transform 1 0 1672 0 1 170
box -8 -3 16 105
use FILL  FILL_1500
timestamp 1681620392
transform 1 0 1680 0 1 170
box -8 -3 16 105
use FILL  FILL_1502
timestamp 1681620392
transform 1 0 1688 0 1 170
box -8 -3 16 105
use FILL  FILL_1504
timestamp 1681620392
transform 1 0 1696 0 1 170
box -8 -3 16 105
use FILL  FILL_1506
timestamp 1681620392
transform 1 0 1704 0 1 170
box -8 -3 16 105
use FILL  FILL_1508
timestamp 1681620392
transform 1 0 1712 0 1 170
box -8 -3 16 105
use FILL  FILL_1510
timestamp 1681620392
transform 1 0 1720 0 1 170
box -8 -3 16 105
use FILL  FILL_1512
timestamp 1681620392
transform 1 0 1728 0 1 170
box -8 -3 16 105
use FILL  FILL_1514
timestamp 1681620392
transform 1 0 1736 0 1 170
box -8 -3 16 105
use FILL  FILL_1516
timestamp 1681620392
transform 1 0 1744 0 1 170
box -8 -3 16 105
use FILL  FILL_1518
timestamp 1681620392
transform 1 0 1752 0 1 170
box -8 -3 16 105
use FILL  FILL_1520
timestamp 1681620392
transform 1 0 1760 0 1 170
box -8 -3 16 105
use FILL  FILL_1522
timestamp 1681620392
transform 1 0 1768 0 1 170
box -8 -3 16 105
use FILL  FILL_1524
timestamp 1681620392
transform 1 0 1776 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_304
timestamp 1681620392
transform 1 0 1784 0 1 170
box -8 -3 104 105
use INVX2  INVX2_373
timestamp 1681620392
transform 1 0 1880 0 1 170
box -9 -3 26 105
use INVX2  INVX2_374
timestamp 1681620392
transform 1 0 1896 0 1 170
box -9 -3 26 105
use M3_M2  M3_M2_4756
timestamp 1681620392
transform 1 0 1940 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_130
timestamp 1681620392
transform -1 0 1952 0 1 170
box -8 -3 46 105
use M3_M2  M3_M2_4757
timestamp 1681620392
transform 1 0 1980 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_131
timestamp 1681620392
transform -1 0 1992 0 1 170
box -8 -3 46 105
use FILL  FILL_1525
timestamp 1681620392
transform 1 0 1992 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_307
timestamp 1681620392
transform 1 0 2000 0 1 170
box -8 -3 104 105
use INVX2  INVX2_376
timestamp 1681620392
transform 1 0 2096 0 1 170
box -9 -3 26 105
use FILL  FILL_1528
timestamp 1681620392
transform 1 0 2112 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_306
timestamp 1681620392
transform 1 0 2120 0 1 170
box -8 -3 34 105
use NAND2X1  NAND2X1_327
timestamp 1681620392
transform -1 0 2176 0 1 170
box -8 -3 32 105
use FILL  FILL_1529
timestamp 1681620392
transform 1 0 2176 0 1 170
box -8 -3 16 105
use FILL  FILL_1541
timestamp 1681620392
transform 1 0 2184 0 1 170
box -8 -3 16 105
use FILL  FILL_1542
timestamp 1681620392
transform 1 0 2192 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_307
timestamp 1681620392
transform 1 0 2200 0 1 170
box -8 -3 34 105
use NAND2X1  NAND2X1_328
timestamp 1681620392
transform -1 0 2256 0 1 170
box -8 -3 32 105
use FILL  FILL_1543
timestamp 1681620392
transform 1 0 2256 0 1 170
box -8 -3 16 105
use FILL  FILL_1544
timestamp 1681620392
transform 1 0 2264 0 1 170
box -8 -3 16 105
use FILL  FILL_1545
timestamp 1681620392
transform 1 0 2272 0 1 170
box -8 -3 16 105
use FILL  FILL_1546
timestamp 1681620392
transform 1 0 2280 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_308
timestamp 1681620392
transform 1 0 2288 0 1 170
box -8 -3 34 105
use M3_M2  M3_M2_4758
timestamp 1681620392
transform 1 0 2348 0 1 175
box -3 -3 3 3
use NAND2X1  NAND2X1_329
timestamp 1681620392
transform -1 0 2344 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_330
timestamp 1681620392
transform -1 0 2368 0 1 170
box -8 -3 32 105
use M3_M2  M3_M2_4759
timestamp 1681620392
transform 1 0 2436 0 1 175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_310
timestamp 1681620392
transform 1 0 2368 0 1 170
box -8 -3 104 105
use FILL  FILL_1548
timestamp 1681620392
transform 1 0 2464 0 1 170
box -8 -3 16 105
use NAND2X1  NAND2X1_331
timestamp 1681620392
transform 1 0 2472 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_332
timestamp 1681620392
transform 1 0 2496 0 1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_309
timestamp 1681620392
transform -1 0 2552 0 1 170
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_311
timestamp 1681620392
transform 1 0 2552 0 1 170
box -8 -3 104 105
use FILL  FILL_1549
timestamp 1681620392
transform 1 0 2648 0 1 170
box -8 -3 16 105
use FILL  FILL_1556
timestamp 1681620392
transform 1 0 2656 0 1 170
box -8 -3 16 105
use FILL  FILL_1558
timestamp 1681620392
transform 1 0 2664 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_312
timestamp 1681620392
transform -1 0 2704 0 1 170
box -8 -3 34 105
use FILL  FILL_1560
timestamp 1681620392
transform 1 0 2704 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_132
timestamp 1681620392
transform 1 0 2712 0 1 170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_314
timestamp 1681620392
transform 1 0 2752 0 1 170
box -8 -3 104 105
use INVX2  INVX2_378
timestamp 1681620392
transform 1 0 2848 0 1 170
box -9 -3 26 105
use FILL  FILL_1562
timestamp 1681620392
transform 1 0 2864 0 1 170
box -8 -3 16 105
use NOR2X1  NOR2X1_115
timestamp 1681620392
transform -1 0 2896 0 1 170
box -8 -3 32 105
use INVX2  INVX2_379
timestamp 1681620392
transform 1 0 2896 0 1 170
box -9 -3 26 105
use OAI21X1  OAI21X1_314
timestamp 1681620392
transform 1 0 2912 0 1 170
box -8 -3 34 105
use INVX2  INVX2_380
timestamp 1681620392
transform -1 0 2960 0 1 170
box -9 -3 26 105
use FILL  FILL_1563
timestamp 1681620392
transform 1 0 2960 0 1 170
box -8 -3 16 105
use FILL  FILL_1564
timestamp 1681620392
transform 1 0 2968 0 1 170
box -8 -3 16 105
use FILL  FILL_1565
timestamp 1681620392
transform 1 0 2976 0 1 170
box -8 -3 16 105
use FILL  FILL_1575
timestamp 1681620392
transform 1 0 2984 0 1 170
box -8 -3 16 105
use FILL  FILL_1577
timestamp 1681620392
transform 1 0 2992 0 1 170
box -8 -3 16 105
use FILL  FILL_1579
timestamp 1681620392
transform 1 0 3000 0 1 170
box -8 -3 16 105
use FILL  FILL_1581
timestamp 1681620392
transform 1 0 3008 0 1 170
box -8 -3 16 105
use Project_Top_VIA0  Project_Top_VIA0_57
timestamp 1681620392
transform 1 0 3043 0 1 170
box -10 -3 10 3
use Project_Top_VIA0  Project_Top_VIA0_58
timestamp 1681620392
transform 1 0 24 0 1 70
box -10 -3 10 3
use FILL  FILL_1435
timestamp 1681620392
transform 1 0 72 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4777
timestamp 1681620392
transform 1 0 92 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_4790
timestamp 1681620392
transform 1 0 140 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5549
timestamp 1681620392
transform 1 0 92 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5604
timestamp 1681620392
transform 1 0 140 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_297
timestamp 1681620392
transform 1 0 80 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_4791
timestamp 1681620392
transform 1 0 188 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5605
timestamp 1681620392
transform 1 0 188 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4845
timestamp 1681620392
transform 1 0 188 0 1 115
box -3 -3 3 3
use FILL  FILL_1436
timestamp 1681620392
transform 1 0 176 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_5606
timestamp 1681620392
transform 1 0 204 0 1 125
box -2 -2 2 2
use INVX2  INVX2_360
timestamp 1681620392
transform 1 0 184 0 -1 170
box -9 -3 26 105
use FILL  FILL_1437
timestamp 1681620392
transform 1 0 200 0 -1 170
box -8 -3 16 105
use FILL  FILL_1438
timestamp 1681620392
transform 1 0 208 0 -1 170
box -8 -3 16 105
use FILL  FILL_1439
timestamp 1681620392
transform 1 0 216 0 -1 170
box -8 -3 16 105
use FILL  FILL_1440
timestamp 1681620392
transform 1 0 224 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_5541
timestamp 1681620392
transform 1 0 252 0 1 145
box -2 -2 2 2
use M3_M2  M3_M2_4792
timestamp 1681620392
transform 1 0 260 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5550
timestamp 1681620392
transform 1 0 260 0 1 135
box -2 -2 2 2
use NOR2X1  NOR2X1_105
timestamp 1681620392
transform -1 0 256 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_4760
timestamp 1681620392
transform 1 0 276 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_5607
timestamp 1681620392
transform 1 0 276 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4846
timestamp 1681620392
transform 1 0 276 0 1 115
box -3 -3 3 3
use NOR2X1  NOR2X1_106
timestamp 1681620392
transform 1 0 256 0 -1 170
box -8 -3 32 105
use M2_M1  M2_M1_5551
timestamp 1681620392
transform 1 0 292 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_4828
timestamp 1681620392
transform 1 0 292 0 1 125
box -3 -3 3 3
use FILL  FILL_1441
timestamp 1681620392
transform 1 0 280 0 -1 170
box -8 -3 16 105
use FILL  FILL_1442
timestamp 1681620392
transform 1 0 288 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4761
timestamp 1681620392
transform 1 0 308 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_5552
timestamp 1681620392
transform 1 0 308 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5608
timestamp 1681620392
transform 1 0 340 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5609
timestamp 1681620392
transform 1 0 388 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4847
timestamp 1681620392
transform 1 0 388 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_298
timestamp 1681620392
transform 1 0 296 0 -1 170
box -8 -3 104 105
use FILL  FILL_1443
timestamp 1681620392
transform 1 0 392 0 -1 170
box -8 -3 16 105
use FILL  FILL_1445
timestamp 1681620392
transform 1 0 400 0 -1 170
box -8 -3 16 105
use FILL  FILL_1446
timestamp 1681620392
transform 1 0 408 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_5542
timestamp 1681620392
transform 1 0 428 0 1 145
box -2 -2 2 2
use FILL  FILL_1447
timestamp 1681620392
transform 1 0 416 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4762
timestamp 1681620392
transform 1 0 460 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_5543
timestamp 1681620392
transform 1 0 444 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_5553
timestamp 1681620392
transform 1 0 452 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5610
timestamp 1681620392
transform 1 0 444 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4829
timestamp 1681620392
transform 1 0 452 0 1 125
box -3 -3 3 3
use NOR2X1  NOR2X1_109
timestamp 1681620392
transform 1 0 424 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_4819
timestamp 1681620392
transform 1 0 484 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_5611
timestamp 1681620392
transform 1 0 468 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5612
timestamp 1681620392
transform 1 0 476 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4848
timestamp 1681620392
transform 1 0 468 0 1 115
box -3 -3 3 3
use NOR2X1  NOR2X1_110
timestamp 1681620392
transform 1 0 448 0 -1 170
box -8 -3 32 105
use FILL  FILL_1449
timestamp 1681620392
transform 1 0 472 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_5554
timestamp 1681620392
transform 1 0 492 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5555
timestamp 1681620392
transform 1 0 500 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_4849
timestamp 1681620392
transform 1 0 500 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_4866
timestamp 1681620392
transform 1 0 492 0 1 105
box -3 -3 3 3
use FILL  FILL_1451
timestamp 1681620392
transform 1 0 480 0 -1 170
box -8 -3 16 105
use FILL  FILL_1453
timestamp 1681620392
transform 1 0 488 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_5544
timestamp 1681620392
transform 1 0 524 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_5613
timestamp 1681620392
transform 1 0 524 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5614
timestamp 1681620392
transform 1 0 532 0 1 125
box -2 -2 2 2
use AOI21X1  AOI21X1_42
timestamp 1681620392
transform 1 0 496 0 -1 170
box -7 -3 39 105
use M3_M2  M3_M2_4793
timestamp 1681620392
transform 1 0 548 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5556
timestamp 1681620392
transform 1 0 540 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5557
timestamp 1681620392
transform 1 0 548 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5615
timestamp 1681620392
transform 1 0 540 0 1 125
box -2 -2 2 2
use INVX2  INVX2_365
timestamp 1681620392
transform -1 0 544 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_4763
timestamp 1681620392
transform 1 0 572 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_5558
timestamp 1681620392
transform 1 0 572 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5616
timestamp 1681620392
transform 1 0 564 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5662
timestamp 1681620392
transform 1 0 572 0 1 115
box -2 -2 2 2
use NAND2X1  NAND2X1_320
timestamp 1681620392
transform 1 0 544 0 -1 170
box -8 -3 32 105
use FILL  FILL_1462
timestamp 1681620392
transform 1 0 568 0 -1 170
box -8 -3 16 105
use FILL  FILL_1463
timestamp 1681620392
transform 1 0 576 0 -1 170
box -8 -3 16 105
use FILL  FILL_1464
timestamp 1681620392
transform 1 0 584 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4850
timestamp 1681620392
transform 1 0 604 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_4794
timestamp 1681620392
transform 1 0 636 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_4820
timestamp 1681620392
transform 1 0 628 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_5559
timestamp 1681620392
transform 1 0 636 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5663
timestamp 1681620392
transform 1 0 612 0 1 115
box -2 -2 2 2
use NAND2X1  NAND2X1_321
timestamp 1681620392
transform 1 0 592 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_4764
timestamp 1681620392
transform 1 0 652 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_5617
timestamp 1681620392
transform 1 0 644 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4830
timestamp 1681620392
transform 1 0 652 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_5545
timestamp 1681620392
transform 1 0 684 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_5618
timestamp 1681620392
transform 1 0 660 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4851
timestamp 1681620392
transform 1 0 644 0 1 115
box -3 -3 3 3
use INVX2  INVX2_366
timestamp 1681620392
transform 1 0 616 0 -1 170
box -9 -3 26 105
use FILL  FILL_1465
timestamp 1681620392
transform 1 0 632 0 -1 170
box -8 -3 16 105
use FILL  FILL_1466
timestamp 1681620392
transform 1 0 640 0 -1 170
box -8 -3 16 105
use AND2X2  AND2X2_31
timestamp 1681620392
transform 1 0 648 0 -1 170
box -8 -3 40 105
use M3_M2  M3_M2_4795
timestamp 1681620392
transform 1 0 708 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5560
timestamp 1681620392
transform 1 0 700 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5561
timestamp 1681620392
transform 1 0 708 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5619
timestamp 1681620392
transform 1 0 700 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4852
timestamp 1681620392
transform 1 0 700 0 1 115
box -3 -3 3 3
use NOR2X1  NOR2X1_111
timestamp 1681620392
transform 1 0 680 0 -1 170
box -8 -3 32 105
use FILL  FILL_1467
timestamp 1681620392
transform 1 0 704 0 -1 170
box -8 -3 16 105
use FILL  FILL_1468
timestamp 1681620392
transform 1 0 712 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4831
timestamp 1681620392
transform 1 0 740 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_5664
timestamp 1681620392
transform 1 0 740 0 1 115
box -2 -2 2 2
use NAND2X1  NAND2X1_322
timestamp 1681620392
transform 1 0 720 0 -1 170
box -8 -3 32 105
use M2_M1  M2_M1_5620
timestamp 1681620392
transform 1 0 756 0 1 125
box -2 -2 2 2
use FILL  FILL_1469
timestamp 1681620392
transform 1 0 744 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4796
timestamp 1681620392
transform 1 0 772 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5546
timestamp 1681620392
transform 1 0 812 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_5562
timestamp 1681620392
transform 1 0 780 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5563
timestamp 1681620392
transform 1 0 796 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_4821
timestamp 1681620392
transform 1 0 804 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_5621
timestamp 1681620392
transform 1 0 772 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5622
timestamp 1681620392
transform 1 0 780 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4867
timestamp 1681620392
transform 1 0 764 0 1 105
box -3 -3 3 3
use FILL  FILL_1470
timestamp 1681620392
transform 1 0 752 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4868
timestamp 1681620392
transform 1 0 780 0 1 105
box -3 -3 3 3
use NAND2X1  NAND2X1_323
timestamp 1681620392
transform -1 0 784 0 -1 170
box -8 -3 32 105
use M2_M1  M2_M1_5623
timestamp 1681620392
transform 1 0 812 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5624
timestamp 1681620392
transform 1 0 820 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4853
timestamp 1681620392
transform 1 0 812 0 1 115
box -3 -3 3 3
use AOI21X1  AOI21X1_43
timestamp 1681620392
transform 1 0 784 0 -1 170
box -7 -3 39 105
use M3_M2  M3_M2_4765
timestamp 1681620392
transform 1 0 836 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_4797
timestamp 1681620392
transform 1 0 828 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5564
timestamp 1681620392
transform 1 0 828 0 1 135
box -2 -2 2 2
use INVX2  INVX2_367
timestamp 1681620392
transform -1 0 832 0 -1 170
box -9 -3 26 105
use M2_M1  M2_M1_5565
timestamp 1681620392
transform 1 0 844 0 1 135
box -2 -2 2 2
use FILL  FILL_1471
timestamp 1681620392
transform 1 0 832 0 -1 170
box -8 -3 16 105
use FILL  FILL_1472
timestamp 1681620392
transform 1 0 840 0 -1 170
box -8 -3 16 105
use FILL  FILL_1473
timestamp 1681620392
transform 1 0 848 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4798
timestamp 1681620392
transform 1 0 884 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5566
timestamp 1681620392
transform 1 0 884 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5625
timestamp 1681620392
transform 1 0 868 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4832
timestamp 1681620392
transform 1 0 884 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_5665
timestamp 1681620392
transform 1 0 884 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_4854
timestamp 1681620392
transform 1 0 892 0 1 115
box -3 -3 3 3
use M2_M1  M2_M1_5683
timestamp 1681620392
transform 1 0 876 0 1 105
box -2 -2 2 2
use INVX2  INVX2_368
timestamp 1681620392
transform 1 0 856 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_4766
timestamp 1681620392
transform 1 0 908 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_5567
timestamp 1681620392
transform 1 0 908 0 1 135
box -2 -2 2 2
use NAND3X1  NAND3X1_124
timestamp 1681620392
transform 1 0 872 0 -1 170
box -8 -3 40 105
use M2_M1  M2_M1_5666
timestamp 1681620392
transform 1 0 916 0 1 115
box -2 -2 2 2
use FILL  FILL_1474
timestamp 1681620392
transform 1 0 904 0 -1 170
box -8 -3 16 105
use FILL  FILL_1475
timestamp 1681620392
transform 1 0 912 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4767
timestamp 1681620392
transform 1 0 940 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_4768
timestamp 1681620392
transform 1 0 956 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_4799
timestamp 1681620392
transform 1 0 940 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5568
timestamp 1681620392
transform 1 0 940 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5569
timestamp 1681620392
transform 1 0 956 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5626
timestamp 1681620392
transform 1 0 932 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4833
timestamp 1681620392
transform 1 0 956 0 1 125
box -3 -3 3 3
use OAI22X1  OAI22X1_129
timestamp 1681620392
transform -1 0 960 0 -1 170
box -8 -3 46 105
use INVX2  INVX2_369
timestamp 1681620392
transform -1 0 976 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_4769
timestamp 1681620392
transform 1 0 996 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_5570
timestamp 1681620392
transform 1 0 988 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_4855
timestamp 1681620392
transform 1 0 988 0 1 115
box -3 -3 3 3
use FILL  FILL_1476
timestamp 1681620392
transform 1 0 976 0 -1 170
box -8 -3 16 105
use FILL  FILL_1477
timestamp 1681620392
transform 1 0 984 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4800
timestamp 1681620392
transform 1 0 1028 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5571
timestamp 1681620392
transform 1 0 1004 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5627
timestamp 1681620392
transform 1 0 1028 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5628
timestamp 1681620392
transform 1 0 1084 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4856
timestamp 1681620392
transform 1 0 1084 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_301
timestamp 1681620392
transform 1 0 992 0 -1 170
box -8 -3 104 105
use FILL  FILL_1478
timestamp 1681620392
transform 1 0 1088 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4801
timestamp 1681620392
transform 1 0 1156 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5572
timestamp 1681620392
transform 1 0 1108 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_4822
timestamp 1681620392
transform 1 0 1188 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_5629
timestamp 1681620392
transform 1 0 1140 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_302
timestamp 1681620392
transform 1 0 1096 0 -1 170
box -8 -3 104 105
use FILL  FILL_1479
timestamp 1681620392
transform 1 0 1192 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4770
timestamp 1681620392
transform 1 0 1212 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_4802
timestamp 1681620392
transform 1 0 1220 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5573
timestamp 1681620392
transform 1 0 1212 0 1 135
box -2 -2 2 2
use FILL  FILL_1480
timestamp 1681620392
transform 1 0 1200 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_5630
timestamp 1681620392
transform 1 0 1220 0 1 125
box -2 -2 2 2
use INVX2  INVX2_370
timestamp 1681620392
transform 1 0 1208 0 -1 170
box -9 -3 26 105
use FILL  FILL_1481
timestamp 1681620392
transform 1 0 1224 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4778
timestamp 1681620392
transform 1 0 1244 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_4779
timestamp 1681620392
transform 1 0 1260 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_4780
timestamp 1681620392
transform 1 0 1332 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_5574
timestamp 1681620392
transform 1 0 1244 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_4823
timestamp 1681620392
transform 1 0 1268 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_5575
timestamp 1681620392
transform 1 0 1332 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5631
timestamp 1681620392
transform 1 0 1268 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5632
timestamp 1681620392
transform 1 0 1332 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5633
timestamp 1681620392
transform 1 0 1340 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_303
timestamp 1681620392
transform 1 0 1232 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_4857
timestamp 1681620392
transform 1 0 1348 0 1 115
box -3 -3 3 3
use INVX2  INVX2_371
timestamp 1681620392
transform 1 0 1328 0 -1 170
box -9 -3 26 105
use FILL  FILL_1482
timestamp 1681620392
transform 1 0 1344 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4771
timestamp 1681620392
transform 1 0 1364 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_5547
timestamp 1681620392
transform 1 0 1364 0 1 145
box -2 -2 2 2
use FILL  FILL_1483
timestamp 1681620392
transform 1 0 1352 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4803
timestamp 1681620392
transform 1 0 1372 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_4781
timestamp 1681620392
transform 1 0 1404 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_5548
timestamp 1681620392
transform 1 0 1380 0 1 145
box -2 -2 2 2
use M3_M2  M3_M2_4804
timestamp 1681620392
transform 1 0 1396 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5576
timestamp 1681620392
transform 1 0 1380 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5577
timestamp 1681620392
transform 1 0 1396 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_4834
timestamp 1681620392
transform 1 0 1380 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_5634
timestamp 1681620392
transform 1 0 1388 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4858
timestamp 1681620392
transform 1 0 1388 0 1 115
box -3 -3 3 3
use NOR2X1  NOR2X1_112
timestamp 1681620392
transform 1 0 1360 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_4782
timestamp 1681620392
transform 1 0 1444 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_4805
timestamp 1681620392
transform 1 0 1460 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5578
timestamp 1681620392
transform 1 0 1420 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5579
timestamp 1681620392
transform 1 0 1444 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5635
timestamp 1681620392
transform 1 0 1404 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4859
timestamp 1681620392
transform 1 0 1404 0 1 115
box -3 -3 3 3
use M2_M1  M2_M1_5667
timestamp 1681620392
transform 1 0 1412 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5684
timestamp 1681620392
transform 1 0 1412 0 1 105
box -2 -2 2 2
use NOR2X1  NOR2X1_113
timestamp 1681620392
transform 1 0 1384 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_4824
timestamp 1681620392
transform 1 0 1452 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_5580
timestamp 1681620392
transform 1 0 1460 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_4825
timestamp 1681620392
transform 1 0 1468 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_5636
timestamp 1681620392
transform 1 0 1444 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4835
timestamp 1681620392
transform 1 0 1460 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_5637
timestamp 1681620392
transform 1 0 1468 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5668
timestamp 1681620392
transform 1 0 1444 0 1 115
box -2 -2 2 2
use NAND3X1  NAND3X1_125
timestamp 1681620392
transform 1 0 1408 0 -1 170
box -8 -3 40 105
use M3_M2  M3_M2_4860
timestamp 1681620392
transform 1 0 1452 0 1 115
box -3 -3 3 3
use M2_M1  M2_M1_5581
timestamp 1681620392
transform 1 0 1484 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_4836
timestamp 1681620392
transform 1 0 1484 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_5669
timestamp 1681620392
transform 1 0 1460 0 1 115
box -2 -2 2 2
use NAND2X1  NAND2X1_324
timestamp 1681620392
transform 1 0 1440 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_4861
timestamp 1681620392
transform 1 0 1476 0 1 115
box -3 -3 3 3
use M2_M1  M2_M1_5670
timestamp 1681620392
transform 1 0 1484 0 1 115
box -2 -2 2 2
use NAND2X1  NAND2X1_325
timestamp 1681620392
transform 1 0 1464 0 -1 170
box -8 -3 32 105
use FILL  FILL_1485
timestamp 1681620392
transform 1 0 1488 0 -1 170
box -8 -3 16 105
use FILL  FILL_1487
timestamp 1681620392
transform 1 0 1496 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_5582
timestamp 1681620392
transform 1 0 1516 0 1 135
box -2 -2 2 2
use FILL  FILL_1488
timestamp 1681620392
transform 1 0 1504 0 -1 170
box -8 -3 16 105
use NAND2X1  NAND2X1_326
timestamp 1681620392
transform 1 0 1512 0 -1 170
box -8 -3 32 105
use FILL  FILL_1489
timestamp 1681620392
transform 1 0 1536 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_5583
timestamp 1681620392
transform 1 0 1564 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_4837
timestamp 1681620392
transform 1 0 1564 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_5671
timestamp 1681620392
transform 1 0 1556 0 1 115
box -2 -2 2 2
use FILL  FILL_1490
timestamp 1681620392
transform 1 0 1544 0 -1 170
box -8 -3 16 105
use FILL  FILL_1491
timestamp 1681620392
transform 1 0 1552 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_5584
timestamp 1681620392
transform 1 0 1588 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_4838
timestamp 1681620392
transform 1 0 1596 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_5638
timestamp 1681620392
transform 1 0 1604 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5672
timestamp 1681620392
transform 1 0 1588 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5673
timestamp 1681620392
transform 1 0 1596 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5674
timestamp 1681620392
transform 1 0 1620 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_4869
timestamp 1681620392
transform 1 0 1588 0 1 105
box -3 -3 3 3
use M2_M1  M2_M1_5685
timestamp 1681620392
transform 1 0 1612 0 1 105
box -2 -2 2 2
use OAI21X1  OAI21X1_305
timestamp 1681620392
transform 1 0 1560 0 -1 170
box -8 -3 34 105
use M3_M2  M3_M2_4870
timestamp 1681620392
transform 1 0 1620 0 1 105
box -3 -3 3 3
use NAND3X1  NAND3X1_128
timestamp 1681620392
transform 1 0 1592 0 -1 170
box -8 -3 40 105
use FILL  FILL_1492
timestamp 1681620392
transform 1 0 1624 0 -1 170
box -8 -3 16 105
use FILL  FILL_1493
timestamp 1681620392
transform 1 0 1632 0 -1 170
box -8 -3 16 105
use FILL  FILL_1495
timestamp 1681620392
transform 1 0 1640 0 -1 170
box -8 -3 16 105
use FILL  FILL_1496
timestamp 1681620392
transform 1 0 1648 0 -1 170
box -8 -3 16 105
use FILL  FILL_1497
timestamp 1681620392
transform 1 0 1656 0 -1 170
box -8 -3 16 105
use FILL  FILL_1498
timestamp 1681620392
transform 1 0 1664 0 -1 170
box -8 -3 16 105
use FILL  FILL_1499
timestamp 1681620392
transform 1 0 1672 0 -1 170
box -8 -3 16 105
use FILL  FILL_1501
timestamp 1681620392
transform 1 0 1680 0 -1 170
box -8 -3 16 105
use FILL  FILL_1503
timestamp 1681620392
transform 1 0 1688 0 -1 170
box -8 -3 16 105
use FILL  FILL_1505
timestamp 1681620392
transform 1 0 1696 0 -1 170
box -8 -3 16 105
use FILL  FILL_1507
timestamp 1681620392
transform 1 0 1704 0 -1 170
box -8 -3 16 105
use FILL  FILL_1509
timestamp 1681620392
transform 1 0 1712 0 -1 170
box -8 -3 16 105
use FILL  FILL_1511
timestamp 1681620392
transform 1 0 1720 0 -1 170
box -8 -3 16 105
use FILL  FILL_1513
timestamp 1681620392
transform 1 0 1728 0 -1 170
box -8 -3 16 105
use FILL  FILL_1515
timestamp 1681620392
transform 1 0 1736 0 -1 170
box -8 -3 16 105
use FILL  FILL_1517
timestamp 1681620392
transform 1 0 1744 0 -1 170
box -8 -3 16 105
use FILL  FILL_1519
timestamp 1681620392
transform 1 0 1752 0 -1 170
box -8 -3 16 105
use FILL  FILL_1521
timestamp 1681620392
transform 1 0 1760 0 -1 170
box -8 -3 16 105
use FILL  FILL_1523
timestamp 1681620392
transform 1 0 1768 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4806
timestamp 1681620392
transform 1 0 1788 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5585
timestamp 1681620392
transform 1 0 1788 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_4807
timestamp 1681620392
transform 1 0 1884 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5586
timestamp 1681620392
transform 1 0 1884 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5639
timestamp 1681620392
transform 1 0 1836 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5640
timestamp 1681620392
transform 1 0 1868 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5641
timestamp 1681620392
transform 1 0 1932 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_305
timestamp 1681620392
transform 1 0 1776 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_306
timestamp 1681620392
transform 1 0 1872 0 -1 170
box -8 -3 104 105
use M2_M1  M2_M1_5642
timestamp 1681620392
transform 1 0 1980 0 1 125
box -2 -2 2 2
use INVX2  INVX2_375
timestamp 1681620392
transform 1 0 1968 0 -1 170
box -9 -3 26 105
use FILL  FILL_1526
timestamp 1681620392
transform 1 0 1984 0 -1 170
box -8 -3 16 105
use FILL  FILL_1527
timestamp 1681620392
transform 1 0 1992 0 -1 170
box -8 -3 16 105
use FILL  FILL_1530
timestamp 1681620392
transform 1 0 2000 0 -1 170
box -8 -3 16 105
use FILL  FILL_1531
timestamp 1681620392
transform 1 0 2008 0 -1 170
box -8 -3 16 105
use FILL  FILL_1532
timestamp 1681620392
transform 1 0 2016 0 -1 170
box -8 -3 16 105
use FILL  FILL_1533
timestamp 1681620392
transform 1 0 2024 0 -1 170
box -8 -3 16 105
use FILL  FILL_1534
timestamp 1681620392
transform 1 0 2032 0 -1 170
box -8 -3 16 105
use FILL  FILL_1535
timestamp 1681620392
transform 1 0 2040 0 -1 170
box -8 -3 16 105
use FILL  FILL_1536
timestamp 1681620392
transform 1 0 2048 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_5643
timestamp 1681620392
transform 1 0 2068 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4862
timestamp 1681620392
transform 1 0 2068 0 1 115
box -3 -3 3 3
use FILL  FILL_1537
timestamp 1681620392
transform 1 0 2056 0 -1 170
box -8 -3 16 105
use FILL  FILL_1538
timestamp 1681620392
transform 1 0 2064 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4808
timestamp 1681620392
transform 1 0 2084 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5587
timestamp 1681620392
transform 1 0 2084 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5644
timestamp 1681620392
transform 1 0 2132 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4826
timestamp 1681620392
transform 1 0 2172 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_5645
timestamp 1681620392
transform 1 0 2172 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_308
timestamp 1681620392
transform 1 0 2072 0 -1 170
box -8 -3 104 105
use FILL  FILL_1539
timestamp 1681620392
transform 1 0 2168 0 -1 170
box -8 -3 16 105
use FILL  FILL_1540
timestamp 1681620392
transform 1 0 2176 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4772
timestamp 1681620392
transform 1 0 2276 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_4809
timestamp 1681620392
transform 1 0 2196 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5588
timestamp 1681620392
transform 1 0 2196 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5589
timestamp 1681620392
transform 1 0 2292 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5646
timestamp 1681620392
transform 1 0 2228 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5647
timestamp 1681620392
transform 1 0 2276 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5648
timestamp 1681620392
transform 1 0 2284 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4863
timestamp 1681620392
transform 1 0 2284 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_309
timestamp 1681620392
transform 1 0 2184 0 -1 170
box -8 -3 104 105
use FILL  FILL_1547
timestamp 1681620392
transform 1 0 2280 0 -1 170
box -8 -3 16 105
use FILL  FILL_1550
timestamp 1681620392
transform 1 0 2288 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4783
timestamp 1681620392
transform 1 0 2348 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_4784
timestamp 1681620392
transform 1 0 2380 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_4810
timestamp 1681620392
transform 1 0 2332 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_4811
timestamp 1681620392
transform 1 0 2372 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5675
timestamp 1681620392
transform 1 0 2324 0 1 115
box -2 -2 2 2
use OAI21X1  OAI21X1_310
timestamp 1681620392
transform 1 0 2296 0 -1 170
box -8 -3 34 105
use M2_M1  M2_M1_5590
timestamp 1681620392
transform 1 0 2332 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5591
timestamp 1681620392
transform 1 0 2348 0 1 135
box -2 -2 2 2
use FILL  FILL_1551
timestamp 1681620392
transform 1 0 2328 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_5649
timestamp 1681620392
transform 1 0 2372 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5592
timestamp 1681620392
transform 1 0 2436 0 1 135
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_312
timestamp 1681620392
transform 1 0 2336 0 -1 170
box -8 -3 104 105
use FILL  FILL_1552
timestamp 1681620392
transform 1 0 2432 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4827
timestamp 1681620392
transform 1 0 2452 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_5593
timestamp 1681620392
transform 1 0 2460 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_4773
timestamp 1681620392
transform 1 0 2492 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_4812
timestamp 1681620392
transform 1 0 2492 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5594
timestamp 1681620392
transform 1 0 2492 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_4839
timestamp 1681620392
transform 1 0 2460 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_5650
timestamp 1681620392
transform 1 0 2468 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5651
timestamp 1681620392
transform 1 0 2476 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4840
timestamp 1681620392
transform 1 0 2484 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_4774
timestamp 1681620392
transform 1 0 2564 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_4785
timestamp 1681620392
transform 1 0 2532 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_4786
timestamp 1681620392
transform 1 0 2564 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_4813
timestamp 1681620392
transform 1 0 2556 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5595
timestamp 1681620392
transform 1 0 2516 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5596
timestamp 1681620392
transform 1 0 2532 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5652
timestamp 1681620392
transform 1 0 2508 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5676
timestamp 1681620392
transform 1 0 2460 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_4864
timestamp 1681620392
transform 1 0 2476 0 1 115
box -3 -3 3 3
use M2_M1  M2_M1_5677
timestamp 1681620392
transform 1 0 2484 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5678
timestamp 1681620392
transform 1 0 2492 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_4871
timestamp 1681620392
transform 1 0 2468 0 1 105
box -3 -3 3 3
use NAND2X1  NAND2X1_333
timestamp 1681620392
transform 1 0 2440 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_4841
timestamp 1681620392
transform 1 0 2516 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_5653
timestamp 1681620392
transform 1 0 2556 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4872
timestamp 1681620392
transform 1 0 2492 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_4873
timestamp 1681620392
transform 1 0 2508 0 1 105
box -3 -3 3 3
use NAND2X1  NAND2X1_334
timestamp 1681620392
transform 1 0 2464 0 -1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_311
timestamp 1681620392
transform -1 0 2520 0 -1 170
box -8 -3 34 105
use M3_M2  M3_M2_4842
timestamp 1681620392
transform 1 0 2620 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_5654
timestamp 1681620392
transform 1 0 2628 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_313
timestamp 1681620392
transform 1 0 2520 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_4865
timestamp 1681620392
transform 1 0 2628 0 1 115
box -3 -3 3 3
use M2_M1  M2_M1_5679
timestamp 1681620392
transform 1 0 2636 0 1 115
box -2 -2 2 2
use INVX2  INVX2_377
timestamp 1681620392
transform 1 0 2616 0 -1 170
box -9 -3 26 105
use FILL  FILL_1553
timestamp 1681620392
transform 1 0 2632 0 -1 170
box -8 -3 16 105
use FILL  FILL_1554
timestamp 1681620392
transform 1 0 2640 0 -1 170
box -8 -3 16 105
use FILL  FILL_1555
timestamp 1681620392
transform 1 0 2648 0 -1 170
box -8 -3 16 105
use FILL  FILL_1557
timestamp 1681620392
transform 1 0 2656 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4814
timestamp 1681620392
transform 1 0 2676 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5597
timestamp 1681620392
transform 1 0 2676 0 1 135
box -2 -2 2 2
use FILL  FILL_1559
timestamp 1681620392
transform 1 0 2664 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_5655
timestamp 1681620392
transform 1 0 2692 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_4874
timestamp 1681620392
transform 1 0 2692 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_4787
timestamp 1681620392
transform 1 0 2708 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_5598
timestamp 1681620392
transform 1 0 2708 0 1 135
box -2 -2 2 2
use OAI21X1  OAI21X1_313
timestamp 1681620392
transform -1 0 2704 0 -1 170
box -8 -3 34 105
use FILL  FILL_1561
timestamp 1681620392
transform 1 0 2704 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4775
timestamp 1681620392
transform 1 0 2724 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_4776
timestamp 1681620392
transform 1 0 2764 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_4788
timestamp 1681620392
transform 1 0 2740 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_4815
timestamp 1681620392
transform 1 0 2748 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5599
timestamp 1681620392
transform 1 0 2724 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5656
timestamp 1681620392
transform 1 0 2748 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5657
timestamp 1681620392
transform 1 0 2812 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_315
timestamp 1681620392
transform 1 0 2712 0 -1 170
box -8 -3 104 105
use FILL  FILL_1566
timestamp 1681620392
transform 1 0 2808 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4789
timestamp 1681620392
transform 1 0 2836 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_4816
timestamp 1681620392
transform 1 0 2828 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5600
timestamp 1681620392
transform 1 0 2828 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5658
timestamp 1681620392
transform 1 0 2836 0 1 125
box -2 -2 2 2
use INVX2  INVX2_381
timestamp 1681620392
transform -1 0 2832 0 -1 170
box -9 -3 26 105
use FILL  FILL_1567
timestamp 1681620392
transform 1 0 2832 0 -1 170
box -8 -3 16 105
use FILL  FILL_1568
timestamp 1681620392
transform 1 0 2840 0 -1 170
box -8 -3 16 105
use FILL  FILL_1569
timestamp 1681620392
transform 1 0 2848 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4843
timestamp 1681620392
transform 1 0 2868 0 1 125
box -3 -3 3 3
use FILL  FILL_1570
timestamp 1681620392
transform 1 0 2856 0 -1 170
box -8 -3 16 105
use FILL  FILL_1571
timestamp 1681620392
transform 1 0 2864 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_4844
timestamp 1681620392
transform 1 0 2892 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_4817
timestamp 1681620392
transform 1 0 2924 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5601
timestamp 1681620392
transform 1 0 2924 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5659
timestamp 1681620392
transform 1 0 2900 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5660
timestamp 1681620392
transform 1 0 2924 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5686
timestamp 1681620392
transform 1 0 2884 0 1 105
box -2 -2 2 2
use FILL  FILL_1572
timestamp 1681620392
transform 1 0 2872 0 -1 170
box -8 -3 16 105
use FILL  FILL_1573
timestamp 1681620392
transform 1 0 2880 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_5680
timestamp 1681620392
transform 1 0 2900 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5681
timestamp 1681620392
transform 1 0 2924 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_4875
timestamp 1681620392
transform 1 0 2924 0 1 105
box -3 -3 3 3
use NAND3X1  NAND3X1_129
timestamp 1681620392
transform 1 0 2888 0 -1 170
box -8 -3 40 105
use M3_M2  M3_M2_4818
timestamp 1681620392
transform 1 0 2940 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_5602
timestamp 1681620392
transform 1 0 2940 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5661
timestamp 1681620392
transform 1 0 2940 0 1 125
box -2 -2 2 2
use NAND2X1  NAND2X1_335
timestamp 1681620392
transform 1 0 2920 0 -1 170
box -8 -3 32 105
use M2_M1  M2_M1_5603
timestamp 1681620392
transform 1 0 2972 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5682
timestamp 1681620392
transform 1 0 2972 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_4876
timestamp 1681620392
transform 1 0 2972 0 1 105
box -3 -3 3 3
use OAI21X1  OAI21X1_315
timestamp 1681620392
transform 1 0 2944 0 -1 170
box -8 -3 34 105
use FILL  FILL_1574
timestamp 1681620392
transform 1 0 2976 0 -1 170
box -8 -3 16 105
use FILL  FILL_1576
timestamp 1681620392
transform 1 0 2984 0 -1 170
box -8 -3 16 105
use FILL  FILL_1578
timestamp 1681620392
transform 1 0 2992 0 -1 170
box -8 -3 16 105
use FILL  FILL_1580
timestamp 1681620392
transform 1 0 3000 0 -1 170
box -8 -3 16 105
use FILL  FILL_1582
timestamp 1681620392
transform 1 0 3008 0 -1 170
box -8 -3 16 105
use Project_Top_VIA0  Project_Top_VIA0_59
timestamp 1681620392
transform 1 0 3067 0 1 70
box -10 -3 10 3
use Project_Top_VIA1  Project_Top_VIA1_4
timestamp 1681620392
transform 1 0 48 0 1 47
box -10 -10 10 10
use Project_Top_VIA1  Project_Top_VIA1_5
timestamp 1681620392
transform 1 0 3043 0 1 47
box -10 -10 10 10
use Project_Top_VIA1  Project_Top_VIA1_6
timestamp 1681620392
transform 1 0 24 0 1 23
box -10 -10 10 10
use Project_Top_VIA1  Project_Top_VIA1_7
timestamp 1681620392
transform 1 0 3067 0 1 23
box -10 -10 10 10
use PadFrame64  PadFrame64_0
timestamp 1681620392
transform 1 0 619 0 1 638
box -2500 -2400 4300 4400
<< labels >>
rlabel metal3 3091 1915 3091 1915 6 in_clka
rlabel metal2 1700 1 1700 1 6 in_clkb
rlabel metal2 604 3038 604 3038 6 in_restart
rlabel metal2 324 3038 324 3038 6 in_start
rlabel metal3 2 2015 2 2015 6 seed[3]
rlabel metal3 2 1925 2 1925 6 seed[2]
rlabel metal3 2 1905 2 1905 6 seed[1]
rlabel metal3 2 1995 2 1995 6 seed[0]
rlabel metal2 476 3038 476 3038 6 P1_no
rlabel metal2 1596 3038 1596 3038 6 P1_decision[2]
rlabel metal2 1580 3038 1580 3038 6 P1_decision[1]
rlabel metal2 1532 3038 1532 3038 6 P1_decision[0]
rlabel metal2 1164 3038 1164 3038 6 num_cards[2]
rlabel metal2 1236 3038 1236 3038 6 num_cards[1]
rlabel metal2 1300 3038 1300 3038 6 num_cards[0]
rlabel metal3 3091 2615 3091 2615 6 P1_out[23]
rlabel metal3 3091 2365 3091 2365 6 P1_out[22]
rlabel metal3 3091 2815 3091 2815 6 P1_out[21]
rlabel metal3 3091 2735 3091 2735 6 P1_out[20]
rlabel metal3 3091 2535 3091 2535 6 P1_out[19]
rlabel metal3 3091 2415 3091 2415 6 P1_out[18]
rlabel metal2 2644 3038 2644 3038 6 P1_out[17]
rlabel metal2 2820 3038 2820 3038 6 P1_out[16]
rlabel metal2 2420 3038 2420 3038 6 P1_out[15]
rlabel metal2 2444 3038 2444 3038 6 P1_out[14]
rlabel metal2 2756 3038 2756 3038 6 P1_out[13]
rlabel metal3 3091 2865 3091 2865 6 P1_out[12]
rlabel metal2 2284 3038 2284 3038 6 P1_out[11]
rlabel metal2 2148 3038 2148 3038 6 P1_out[10]
rlabel metal2 1924 3038 1924 3038 6 P1_out[9]
rlabel metal2 2028 3038 2028 3038 6 P1_out[8]
rlabel metal2 2100 3038 2100 3038 6 P1_out[7]
rlabel metal2 2268 3038 2268 3038 6 P1_out[6]
rlabel metal2 1852 3038 1852 3038 6 P1_out[5]
rlabel metal2 1500 3038 1500 3038 6 P1_out[4]
rlabel metal2 1476 3038 1476 3038 6 P1_out[3]
rlabel metal2 1460 3038 1460 3038 6 P1_out[2]
rlabel metal2 1516 3038 1516 3038 6 P1_out[1]
rlabel metal2 1380 3038 1380 3038 6 P1_out[0]
rlabel metal3 3091 2165 3091 2165 6 max_card[5]
rlabel metal3 3091 2015 3091 2015 6 max_card[4]
rlabel metal3 3091 1935 3091 1935 6 max_card[3]
rlabel metal3 3091 2265 3091 2265 6 max_card[2]
rlabel metal3 3091 2185 3091 2185 6 max_card[1]
rlabel metal3 3091 2145 3091 2145 6 max_card[0]
rlabel metal2 836 3038 836 3038 6 P2_num_cards[2]
rlabel metal2 860 3038 860 3038 6 P2_num_cards[1]
rlabel metal2 748 3038 748 3038 6 P2_num_cards[0]
rlabel metal3 2 2365 2 2365 6 winner[1]
rlabel metal3 2 2295 2 2295 6 winner[0]
rlabel metal1 38 167 38 167 6 gnd
rlabel metal1 14 67 14 67 6 vdd
rlabel metal1 -130 -1471 -130 -1471 2 p_in_clkb
rlabel metal1 -1587 887 -1587 887 4 GND!
rlabel metal1 -1586 1188 -1586 1188 4 p_P1_no
rlabel metal1 -1589 1486 -1589 1486 4 p_in_restart
rlabel metal1 -1583 2691 -1583 2691 4 GND!
rlabel metal1 3169 4742 3169 4742 6 Vdd!
rlabel metal1 1069 4742 1069 4742 6 Vdd!
rlabel metal1 4624 2385 4624 2385 6 GND!
rlabel metal1 4624 586 4624 586 6 GND!
rlabel metal1 2569 -1476 2569 -1476 8 p_in_clka
rlabel metal1 468 -1468 468 -1468 8 Vdd!
rlabel metal1 2269 -1473 2269 -1473 8 Vdd!
rlabel metal1 -431 -1468 -431 -1468 2 p_seed[1]
rlabel metal1 -731 -1466 -731 -1466 2 p_seed[2]
rlabel metal1 -1586 -611 -1586 -611 2 p_seed[0]
rlabel metal1 -1590 -314 -1590 -314 2 p_seed[3]
rlabel metal1 -1588 -11 -1588 -11 2 p_winner[0]
rlabel metal1 -1586 287 -1586 287 4 p_winner[1]
rlabel metal1 -1589 586 -1589 586 4 p_in_start
rlabel metal1 -1592 1790 -1592 1790 4 p_P2_num_cards[0]
rlabel metal1 -1590 2088 -1590 2088 4 p_P2_num_cards[2]
rlabel metal1 -1587 2389 -1587 2389 4 p_P2_num_cards[1]
rlabel metal1 -1587 2984 -1587 2984 4 p_num_cards[2]
rlabel metal1 -1590 3284 -1590 3284 4 p_num_cards[1]
rlabel metal1 -1593 3586 -1593 3586 4 p_num_cards[0]
rlabel metal1 -1590 3886 -1590 3886 4 p_P1_out[0]
rlabel metal1 -731 4745 -731 4745 4 p_P1_out[2]
rlabel metal1 -428 4748 -428 4748 4 p_P1_out[3]
rlabel metal1 -132 4745 -132 4745 4 p_P1_out[4]
rlabel metal1 168 4744 168 4744 6 p_P1_out[1]
rlabel metal1 466 4747 466 4747 6 p_P1_decision[0]
rlabel metal1 773 4746 773 4746 6 p_P1_decision[1]
rlabel metal1 1370 4747 1370 4747 6 p_P1_decision[2]
rlabel metal1 1669 4745 1669 4745 6 p_P1_out[5]
rlabel metal1 1969 4744 1969 4744 6 p_P1_out[9]
rlabel metal1 2273 4741 2273 4741 6 p_P1_out[8]
rlabel metal1 2569 4749 2569 4749 6 p_P1_out[7]
rlabel metal1 2870 4745 2870 4745 6 p_P1_out[10]
rlabel metal1 3471 4743 3471 4743 6 p_P1_out[6]
rlabel metal1 3769 4747 3769 4747 6 p_P1_out[11]
rlabel metal1 4624 3884 4624 3884 6 p_P1_out[15]
rlabel metal1 4628 2989 4628 2989 6 p_P1_out[13]
rlabel metal1 4625 3281 4625 3281 6 p_P1_out[17]
rlabel metal1 4620 3584 4620 3584 6 p_P1_out[14]
rlabel metal1 4626 2687 4626 2687 6 p_P1_out[16]
rlabel metal1 4626 2087 4626 2087 6 p_P1_out[12]
rlabel metal1 4627 1788 4627 1788 6 p_P1_out[21]
rlabel metal1 4630 1489 4630 1489 6 p_P1_out[20]
rlabel metal1 4627 1185 4627 1185 6 p_P1_out[23]
rlabel metal1 4624 886 4624 886 6 p_P1_out[19]
rlabel metal1 4629 284 4629 284 6 p_P1_out[18]
rlabel metal1 4631 -13 4631 -13 8 p_P1_out[22]
rlabel metal1 4626 -312 4626 -312 8 p_max_card[2]
rlabel metal1 4627 -616 4627 -616 8 p_max_card[1]
rlabel metal1 3769 -1470 3769 -1470 8 p_max_card[5]
rlabel metal1 3470 -1472 3470 -1472 8 p_max_card[0]
rlabel metal1 3169 -1475 3169 -1475 8 p_max_card[4]
rlabel metal1 2869 -1474 2869 -1474 8 p_max_card[3]
<< end >>
