magic
tech scmos
timestamp 1681620392
<< nwell >>
rect -5 48 28 105
<< ntransistor >>
rect 7 6 9 16
rect 15 6 17 26
<< ptransistor >>
rect 7 74 9 94
rect 15 54 17 94
<< ndiffusion >>
rect 10 16 15 26
rect 2 6 7 16
rect 9 6 15 16
rect 17 6 22 26
<< pdiffusion >>
rect 2 74 7 94
rect 9 74 15 94
rect 10 54 15 74
rect 17 54 22 94
<< psubstratepdiff >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratendiff >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 7 57 9 74
rect 6 55 9 57
rect 6 43 8 55
rect 15 51 17 54
rect 12 47 17 51
rect 2 41 8 43
rect 2 39 9 41
rect 7 16 9 39
rect 15 26 17 47
rect 7 4 9 6
rect 15 4 17 6
<< genericcontact >>
rect -1 99 1 101
rect 15 99 17 101
rect 3 90 5 92
rect 11 91 13 93
rect 19 90 21 92
rect 3 85 5 87
rect 11 86 13 88
rect 19 85 21 87
rect 3 80 5 82
rect 11 81 13 83
rect 19 80 21 82
rect 3 75 5 77
rect 11 76 13 78
rect 19 75 21 77
rect 11 71 13 73
rect 19 70 21 72
rect 11 66 13 68
rect 19 65 21 67
rect 11 61 13 63
rect 19 60 21 62
rect 19 55 21 57
rect 13 48 15 50
rect 3 40 5 42
rect 11 22 13 24
rect 19 22 21 24
rect 11 17 13 19
rect 19 17 21 19
rect 3 12 5 14
rect 11 12 13 14
rect 19 12 21 14
rect 3 7 5 9
rect 11 7 13 9
rect 19 7 21 9
rect -1 -1 1 1
rect 15 -1 17 1
<< metal1 >>
rect -2 97 26 103
rect 2 57 6 94
rect 10 60 14 97
rect 2 54 13 57
rect 18 54 22 94
rect 10 51 13 54
rect 10 47 16 51
rect 2 39 6 47
rect 10 32 13 47
rect 19 43 22 54
rect 2 29 13 32
rect 2 6 6 29
rect 10 3 14 26
rect 18 6 22 43
rect -2 -3 26 3
<< m1p >>
rect 2 43 6 47
rect 18 33 22 37
<< labels >>
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 4 0 4 0 8 gnd
rlabel metal1 4 45 4 45 6 A
rlabel metal1 20 35 20 35 6 Y
<< end >>
